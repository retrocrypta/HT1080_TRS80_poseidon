library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0e0c287",
    12 => x"86c0c84e",
    13 => x"49f0e0c2",
    14 => x"48f0cec2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c8dd",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"c44a711e",
    47 => x"c1484966",
    48 => x"58a6c888",
    49 => x"d6029971",
    50 => x"48d4ff87",
    51 => x"6878ffc3",
    52 => x"4966c452",
    53 => x"c888c148",
    54 => x"997158a6",
    55 => x"2687ea05",
    56 => x"1e731e4f",
    57 => x"c34bd4ff",
    58 => x"4a6b7bff",
    59 => x"6b7bffc3",
    60 => x"7232c849",
    61 => x"7bffc3b1",
    62 => x"31c84a6b",
    63 => x"ffc3b271",
    64 => x"c8496b7b",
    65 => x"71b17232",
    66 => x"2687c448",
    67 => x"264c264d",
    68 => x"0e4f264b",
    69 => x"5d5c5b5e",
    70 => x"ff4a710e",
    71 => x"49724cd4",
    72 => x"7199ffc3",
    73 => x"f0cec27c",
    74 => x"87c805bf",
    75 => x"c94866d0",
    76 => x"58a6d430",
    77 => x"d84966d0",
    78 => x"99ffc329",
    79 => x"66d07c71",
    80 => x"c329d049",
    81 => x"7c7199ff",
    82 => x"c84966d0",
    83 => x"99ffc329",
    84 => x"66d07c71",
    85 => x"99ffc349",
    86 => x"49727c71",
    87 => x"ffc329d0",
    88 => x"6c7c7199",
    89 => x"fff0c94b",
    90 => x"abffc34d",
    91 => x"c387d005",
    92 => x"4b6c7cff",
    93 => x"c6028dc1",
    94 => x"abffc387",
    95 => x"7387f002",
    96 => x"87c7fe48",
    97 => x"ff49c01e",
    98 => x"ffc348d4",
    99 => x"c381c178",
   100 => x"04a9b7c8",
   101 => x"4f2687f1",
   102 => x"e71e731e",
   103 => x"dff8c487",
   104 => x"c01ec04b",
   105 => x"f7c1f0ff",
   106 => x"87e7fd49",
   107 => x"a8c186c4",
   108 => x"87eac005",
   109 => x"c348d4ff",
   110 => x"c0c178ff",
   111 => x"c0c0c0c0",
   112 => x"f0e1c01e",
   113 => x"fd49e9c1",
   114 => x"86c487c9",
   115 => x"ca059870",
   116 => x"48d4ff87",
   117 => x"c178ffc3",
   118 => x"fe87cb48",
   119 => x"8bc187e6",
   120 => x"87fdfe05",
   121 => x"e6fc48c0",
   122 => x"1e731e87",
   123 => x"c348d4ff",
   124 => x"4bd378ff",
   125 => x"ffc01ec0",
   126 => x"49c1c1f0",
   127 => x"c487d4fc",
   128 => x"05987086",
   129 => x"d4ff87ca",
   130 => x"78ffc348",
   131 => x"87cb48c1",
   132 => x"c187f1fd",
   133 => x"dbff058b",
   134 => x"fb48c087",
   135 => x"5e0e87f1",
   136 => x"ff0e5c5b",
   137 => x"dbfd4cd4",
   138 => x"1eeac687",
   139 => x"c1f0e1c0",
   140 => x"defb49c8",
   141 => x"c186c487",
   142 => x"87c802a8",
   143 => x"c087eafe",
   144 => x"87e2c148",
   145 => x"7087dafa",
   146 => x"ffffcf49",
   147 => x"a9eac699",
   148 => x"fe87c802",
   149 => x"48c087d3",
   150 => x"c387cbc1",
   151 => x"f1c07cff",
   152 => x"87f4fc4b",
   153 => x"c0029870",
   154 => x"1ec087eb",
   155 => x"c1f0ffc0",
   156 => x"defa49fa",
   157 => x"7086c487",
   158 => x"87d90598",
   159 => x"6c7cffc3",
   160 => x"7cffc349",
   161 => x"c17c7c7c",
   162 => x"c40299c0",
   163 => x"d548c187",
   164 => x"d148c087",
   165 => x"05abc287",
   166 => x"48c087c4",
   167 => x"8bc187c8",
   168 => x"87fdfe05",
   169 => x"e4f948c0",
   170 => x"1e731e87",
   171 => x"48f0cec2",
   172 => x"4bc778c1",
   173 => x"c248d0ff",
   174 => x"87c8fb78",
   175 => x"c348d0ff",
   176 => x"c01ec078",
   177 => x"c0c1d0e5",
   178 => x"87c7f949",
   179 => x"a8c186c4",
   180 => x"4b87c105",
   181 => x"c505abc2",
   182 => x"c048c087",
   183 => x"8bc187f9",
   184 => x"87d0ff05",
   185 => x"c287f7fc",
   186 => x"7058f4ce",
   187 => x"87cd0598",
   188 => x"ffc01ec1",
   189 => x"49d0c1f0",
   190 => x"c487d8f8",
   191 => x"48d4ff86",
   192 => x"c278ffc3",
   193 => x"cec287fc",
   194 => x"d0ff58f8",
   195 => x"ff78c248",
   196 => x"ffc348d4",
   197 => x"f748c178",
   198 => x"5e0e87f5",
   199 => x"0e5d5c5b",
   200 => x"4cc04b71",
   201 => x"dfcdeec5",
   202 => x"48d4ff4a",
   203 => x"6878ffc3",
   204 => x"a9fec349",
   205 => x"87fdc005",
   206 => x"9b734d70",
   207 => x"d087cc02",
   208 => x"49731e66",
   209 => x"c487f1f5",
   210 => x"ff87d686",
   211 => x"d1c448d0",
   212 => x"7dffc378",
   213 => x"c14866d0",
   214 => x"58a6d488",
   215 => x"f0059870",
   216 => x"48d4ff87",
   217 => x"7878ffc3",
   218 => x"c5059b73",
   219 => x"48d0ff87",
   220 => x"4ac178d0",
   221 => x"058ac14c",
   222 => x"7487eefe",
   223 => x"87cbf648",
   224 => x"711e731e",
   225 => x"ff4bc04a",
   226 => x"ffc348d4",
   227 => x"48d0ff78",
   228 => x"ff78c3c4",
   229 => x"ffc348d4",
   230 => x"c01e7278",
   231 => x"d1c1f0ff",
   232 => x"87eff549",
   233 => x"987086c4",
   234 => x"c887d205",
   235 => x"66cc1ec0",
   236 => x"87e6fd49",
   237 => x"4b7086c4",
   238 => x"c248d0ff",
   239 => x"f5487378",
   240 => x"5e0e87cd",
   241 => x"0e5d5c5b",
   242 => x"ffc01ec0",
   243 => x"49c9c1f0",
   244 => x"d287c0f5",
   245 => x"f8cec21e",
   246 => x"87fefc49",
   247 => x"4cc086c8",
   248 => x"b7d284c1",
   249 => x"87f804ac",
   250 => x"97f8cec2",
   251 => x"c0c349bf",
   252 => x"a9c0c199",
   253 => x"87e7c005",
   254 => x"97ffcec2",
   255 => x"31d049bf",
   256 => x"97c0cfc2",
   257 => x"32c84abf",
   258 => x"cfc2b172",
   259 => x"4abf97c1",
   260 => x"cf4c71b1",
   261 => x"9cffffff",
   262 => x"34ca84c1",
   263 => x"c287e7c1",
   264 => x"bf97c1cf",
   265 => x"c631c149",
   266 => x"c2cfc299",
   267 => x"c74abf97",
   268 => x"b1722ab7",
   269 => x"97fdcec2",
   270 => x"cf4d4abf",
   271 => x"fecec29d",
   272 => x"c34abf97",
   273 => x"c232ca9a",
   274 => x"bf97ffce",
   275 => x"7333c24b",
   276 => x"c0cfc2b2",
   277 => x"c34bbf97",
   278 => x"b7c69bc0",
   279 => x"c2b2732b",
   280 => x"7148c181",
   281 => x"c1497030",
   282 => x"70307548",
   283 => x"c14c724d",
   284 => x"c8947184",
   285 => x"06adb7c0",
   286 => x"34c187cc",
   287 => x"c0c82db7",
   288 => x"ff01adb7",
   289 => x"487487f4",
   290 => x"0e87c0f2",
   291 => x"5d5c5b5e",
   292 => x"c286f80e",
   293 => x"c048ded7",
   294 => x"d6cfc278",
   295 => x"fb49c01e",
   296 => x"86c487de",
   297 => x"c5059870",
   298 => x"c948c087",
   299 => x"4dc087ce",
   300 => x"edc07ec1",
   301 => x"c249bff3",
   302 => x"714accd0",
   303 => x"e9ee4bc8",
   304 => x"05987087",
   305 => x"7ec087c2",
   306 => x"bfefedc0",
   307 => x"e8d0c249",
   308 => x"4bc8714a",
   309 => x"7087d3ee",
   310 => x"87c20598",
   311 => x"026e7ec0",
   312 => x"c287fdc0",
   313 => x"4dbfdcd6",
   314 => x"9fd4d7c2",
   315 => x"c5487ebf",
   316 => x"05a8ead6",
   317 => x"d6c287c7",
   318 => x"ce4dbfdc",
   319 => x"ca486e87",
   320 => x"02a8d5e9",
   321 => x"48c087c5",
   322 => x"c287f1c7",
   323 => x"751ed6cf",
   324 => x"87ecf949",
   325 => x"987086c4",
   326 => x"c087c505",
   327 => x"87dcc748",
   328 => x"bfefedc0",
   329 => x"e8d0c249",
   330 => x"4bc8714a",
   331 => x"7087fbec",
   332 => x"87c80598",
   333 => x"48ded7c2",
   334 => x"87da78c1",
   335 => x"bff3edc0",
   336 => x"ccd0c249",
   337 => x"4bc8714a",
   338 => x"7087dfec",
   339 => x"c5c00298",
   340 => x"c648c087",
   341 => x"d7c287e6",
   342 => x"49bf97d4",
   343 => x"05a9d5c1",
   344 => x"c287cdc0",
   345 => x"bf97d5d7",
   346 => x"a9eac249",
   347 => x"87c5c002",
   348 => x"c7c648c0",
   349 => x"d6cfc287",
   350 => x"487ebf97",
   351 => x"02a8e9c3",
   352 => x"6e87cec0",
   353 => x"a8ebc348",
   354 => x"87c5c002",
   355 => x"ebc548c0",
   356 => x"e1cfc287",
   357 => x"9949bf97",
   358 => x"87ccc005",
   359 => x"97e2cfc2",
   360 => x"a9c249bf",
   361 => x"87c5c002",
   362 => x"cfc548c0",
   363 => x"e3cfc287",
   364 => x"c248bf97",
   365 => x"7058dad7",
   366 => x"88c1484c",
   367 => x"58ded7c2",
   368 => x"97e4cfc2",
   369 => x"817549bf",
   370 => x"97e5cfc2",
   371 => x"32c84abf",
   372 => x"c27ea172",
   373 => x"6e48ebdb",
   374 => x"e6cfc278",
   375 => x"c848bf97",
   376 => x"d7c258a6",
   377 => x"c202bfde",
   378 => x"edc087d4",
   379 => x"c249bfef",
   380 => x"714ae8d0",
   381 => x"f1e94bc8",
   382 => x"02987087",
   383 => x"c087c5c0",
   384 => x"87f8c348",
   385 => x"bfd6d7c2",
   386 => x"ffdbc24c",
   387 => x"fbcfc25c",
   388 => x"c849bf97",
   389 => x"facfc231",
   390 => x"a14abf97",
   391 => x"fccfc249",
   392 => x"d04abf97",
   393 => x"49a17232",
   394 => x"97fdcfc2",
   395 => x"32d84abf",
   396 => x"c449a172",
   397 => x"dbc29166",
   398 => x"c281bfeb",
   399 => x"c259f3db",
   400 => x"bf97c3d0",
   401 => x"c232c84a",
   402 => x"bf97c2d0",
   403 => x"c24aa24b",
   404 => x"bf97c4d0",
   405 => x"7333d04b",
   406 => x"d0c24aa2",
   407 => x"4bbf97c5",
   408 => x"33d89bcf",
   409 => x"c24aa273",
   410 => x"c25af7db",
   411 => x"4abff3db",
   412 => x"92748ac2",
   413 => x"48f7dbc2",
   414 => x"c178a172",
   415 => x"cfc287ca",
   416 => x"49bf97e8",
   417 => x"cfc231c8",
   418 => x"4abf97e7",
   419 => x"d7c249a1",
   420 => x"d7c259e6",
   421 => x"c549bfe2",
   422 => x"81ffc731",
   423 => x"dbc229c9",
   424 => x"cfc259ff",
   425 => x"4abf97ed",
   426 => x"cfc232c8",
   427 => x"4bbf97ec",
   428 => x"66c44aa2",
   429 => x"c2826e92",
   430 => x"c25afbdb",
   431 => x"c048f3db",
   432 => x"efdbc278",
   433 => x"78a17248",
   434 => x"48ffdbc2",
   435 => x"bff3dbc2",
   436 => x"c3dcc278",
   437 => x"f7dbc248",
   438 => x"d7c278bf",
   439 => x"c002bfde",
   440 => x"487487c9",
   441 => x"7e7030c4",
   442 => x"c287c9c0",
   443 => x"48bffbdb",
   444 => x"7e7030c4",
   445 => x"48e2d7c2",
   446 => x"48c1786e",
   447 => x"4d268ef8",
   448 => x"4b264c26",
   449 => x"5e0e4f26",
   450 => x"0e5d5c5b",
   451 => x"d7c24a71",
   452 => x"cb02bfde",
   453 => x"c74b7287",
   454 => x"c14c722b",
   455 => x"87c99cff",
   456 => x"2bc84b72",
   457 => x"ffc34c72",
   458 => x"ebdbc29c",
   459 => x"edc083bf",
   460 => x"02abbfeb",
   461 => x"edc087d9",
   462 => x"cfc25bef",
   463 => x"49731ed6",
   464 => x"c487fdf0",
   465 => x"05987086",
   466 => x"48c087c5",
   467 => x"c287e6c0",
   468 => x"02bfded7",
   469 => x"497487d2",
   470 => x"cfc291c4",
   471 => x"4d6981d6",
   472 => x"ffffffcf",
   473 => x"87cb9dff",
   474 => x"91c24974",
   475 => x"81d6cfc2",
   476 => x"754d699f",
   477 => x"87c6fe48",
   478 => x"5c5b5e0e",
   479 => x"86f80e5d",
   480 => x"059c4c71",
   481 => x"48c087c5",
   482 => x"c887c1c3",
   483 => x"486e7ea4",
   484 => x"66d878c0",
   485 => x"d887c702",
   486 => x"05bf9766",
   487 => x"48c087c5",
   488 => x"c087e9c2",
   489 => x"c749c11e",
   490 => x"86c487e6",
   491 => x"029d4d70",
   492 => x"c287c2c1",
   493 => x"d84ae6d7",
   494 => x"d2e24966",
   495 => x"02987087",
   496 => x"7587f2c0",
   497 => x"4966d84a",
   498 => x"f7e24bcb",
   499 => x"02987087",
   500 => x"c087e2c0",
   501 => x"029d751e",
   502 => x"a6c887c7",
   503 => x"c578c048",
   504 => x"48a6c887",
   505 => x"66c878c1",
   506 => x"87e4c649",
   507 => x"4d7086c4",
   508 => x"fefe059d",
   509 => x"029d7587",
   510 => x"dc87cfc1",
   511 => x"486e49a5",
   512 => x"a5da7869",
   513 => x"48a6c449",
   514 => x"9f78a4c4",
   515 => x"66c44869",
   516 => x"d7c27808",
   517 => x"d202bfde",
   518 => x"49a5d487",
   519 => x"c049699f",
   520 => x"7199ffff",
   521 => x"7030d048",
   522 => x"c087c27e",
   523 => x"48496e7e",
   524 => x"80bf66c4",
   525 => x"780866c4",
   526 => x"a4cc7cc0",
   527 => x"bf66c449",
   528 => x"49a4d079",
   529 => x"48c179c0",
   530 => x"48c087c2",
   531 => x"edfa8ef8",
   532 => x"5b5e0e87",
   533 => x"710e5d5c",
   534 => x"c1029c4c",
   535 => x"a4c887ca",
   536 => x"c1026949",
   537 => x"66d087c2",
   538 => x"82496c4a",
   539 => x"d05aa6d4",
   540 => x"c2b94d66",
   541 => x"4abfdad7",
   542 => x"9972baff",
   543 => x"c0029971",
   544 => x"a4c487e4",
   545 => x"f9496b4b",
   546 => x"7b7087fc",
   547 => x"bfd6d7c2",
   548 => x"71816c49",
   549 => x"c2b9757c",
   550 => x"4abfdad7",
   551 => x"9972baff",
   552 => x"ff059971",
   553 => x"7c7587dc",
   554 => x"1e87d3f9",
   555 => x"4b711e73",
   556 => x"87c7029b",
   557 => x"6949a3c8",
   558 => x"c087c505",
   559 => x"87f7c048",
   560 => x"bfefdbc2",
   561 => x"49a3c44a",
   562 => x"89c24969",
   563 => x"bfd6d7c2",
   564 => x"4aa27191",
   565 => x"bfdad7c2",
   566 => x"71996b49",
   567 => x"edc04aa2",
   568 => x"66c85aef",
   569 => x"ea49721e",
   570 => x"86c487d6",
   571 => x"c4059870",
   572 => x"c248c087",
   573 => x"f848c187",
   574 => x"731e87c8",
   575 => x"9b4b711e",
   576 => x"87e4c002",
   577 => x"5bc3dcc2",
   578 => x"8ac24a73",
   579 => x"bfd6d7c2",
   580 => x"dbc29249",
   581 => x"7248bfef",
   582 => x"c7dcc280",
   583 => x"c4487158",
   584 => x"e6d7c230",
   585 => x"87edc058",
   586 => x"48ffdbc2",
   587 => x"bff3dbc2",
   588 => x"c3dcc278",
   589 => x"f7dbc248",
   590 => x"d7c278bf",
   591 => x"c902bfde",
   592 => x"d6d7c287",
   593 => x"31c449bf",
   594 => x"dbc287c7",
   595 => x"c449bffb",
   596 => x"e6d7c231",
   597 => x"87eaf659",
   598 => x"5c5b5e0e",
   599 => x"c04a710e",
   600 => x"029a724b",
   601 => x"da87e1c0",
   602 => x"699f49a2",
   603 => x"ded7c24b",
   604 => x"87cf02bf",
   605 => x"9f49a2d4",
   606 => x"c04c4969",
   607 => x"d09cffff",
   608 => x"c087c234",
   609 => x"b349744c",
   610 => x"edfd4973",
   611 => x"87f0f587",
   612 => x"5c5b5e0e",
   613 => x"86f40e5d",
   614 => x"7ec04a71",
   615 => x"d8029a72",
   616 => x"d2cfc287",
   617 => x"c278c048",
   618 => x"c248cacf",
   619 => x"78bfc3dc",
   620 => x"48cecfc2",
   621 => x"bfffdbc2",
   622 => x"f3d7c278",
   623 => x"c250c048",
   624 => x"49bfe2d7",
   625 => x"bfd2cfc2",
   626 => x"03aa714a",
   627 => x"7287c9c4",
   628 => x"0599cf49",
   629 => x"c087e9c0",
   630 => x"c248ebed",
   631 => x"78bfcacf",
   632 => x"1ed6cfc2",
   633 => x"bfcacfc2",
   634 => x"cacfc249",
   635 => x"78a1c148",
   636 => x"87cce671",
   637 => x"edc086c4",
   638 => x"cfc248e7",
   639 => x"87cc78d6",
   640 => x"bfe7edc0",
   641 => x"80e0c048",
   642 => x"58ebedc0",
   643 => x"bfd2cfc2",
   644 => x"c280c148",
   645 => x"2758d6cf",
   646 => x"00000b67",
   647 => x"4dbf97bf",
   648 => x"e3c2029d",
   649 => x"ade5c387",
   650 => x"87dcc202",
   651 => x"bfe7edc0",
   652 => x"49a3cb4b",
   653 => x"accf4c11",
   654 => x"87d2c105",
   655 => x"99df4975",
   656 => x"91cd89c1",
   657 => x"81e6d7c2",
   658 => x"124aa3c1",
   659 => x"4aa3c351",
   660 => x"a3c55112",
   661 => x"c751124a",
   662 => x"51124aa3",
   663 => x"124aa3c9",
   664 => x"4aa3ce51",
   665 => x"a3d05112",
   666 => x"d251124a",
   667 => x"51124aa3",
   668 => x"124aa3d4",
   669 => x"4aa3d651",
   670 => x"a3d85112",
   671 => x"dc51124a",
   672 => x"51124aa3",
   673 => x"124aa3de",
   674 => x"c07ec151",
   675 => x"497487fa",
   676 => x"c00599c8",
   677 => x"497487eb",
   678 => x"d10599d0",
   679 => x"0266dc87",
   680 => x"7387cbc0",
   681 => x"0f66dc49",
   682 => x"c0029870",
   683 => x"056e87d3",
   684 => x"c287c6c0",
   685 => x"c048e6d7",
   686 => x"e7edc050",
   687 => x"e1c248bf",
   688 => x"f3d7c287",
   689 => x"7e50c048",
   690 => x"bfe2d7c2",
   691 => x"d2cfc249",
   692 => x"aa714abf",
   693 => x"87f7fb04",
   694 => x"bfc3dcc2",
   695 => x"87c8c005",
   696 => x"bfded7c2",
   697 => x"87f8c102",
   698 => x"bfcecfc2",
   699 => x"87d6f049",
   700 => x"cfc24970",
   701 => x"a6c459d2",
   702 => x"cecfc248",
   703 => x"d7c278bf",
   704 => x"c002bfde",
   705 => x"66c487d8",
   706 => x"ffffcf49",
   707 => x"a999f8ff",
   708 => x"87c5c002",
   709 => x"e1c04cc0",
   710 => x"c04cc187",
   711 => x"66c487dc",
   712 => x"f8ffcf49",
   713 => x"c002a999",
   714 => x"a6c887c8",
   715 => x"c078c048",
   716 => x"a6c887c5",
   717 => x"c878c148",
   718 => x"9c744c66",
   719 => x"87e0c005",
   720 => x"c24966c4",
   721 => x"d6d7c289",
   722 => x"c2914abf",
   723 => x"4abfefdb",
   724 => x"48cacfc2",
   725 => x"c278a172",
   726 => x"c048d2cf",
   727 => x"87dff978",
   728 => x"8ef448c0",
   729 => x"0087d7ee",
   730 => x"ff000000",
   731 => x"77ffffff",
   732 => x"8000000b",
   733 => x"4600000b",
   734 => x"32335441",
   735 => x"00202020",
   736 => x"31544146",
   737 => x"20202036",
   738 => x"d4ff1e00",
   739 => x"78ffc348",
   740 => x"4f264868",
   741 => x"48d4ff1e",
   742 => x"ff78ffc3",
   743 => x"e1c048d0",
   744 => x"48d4ff78",
   745 => x"dcc278d4",
   746 => x"d4ff48c7",
   747 => x"4f2650bf",
   748 => x"48d0ff1e",
   749 => x"2678e0c0",
   750 => x"ccff1e4f",
   751 => x"99497087",
   752 => x"c087c602",
   753 => x"f105a9fb",
   754 => x"26487187",
   755 => x"5b5e0e4f",
   756 => x"4b710e5c",
   757 => x"f0fe4cc0",
   758 => x"99497087",
   759 => x"87f9c002",
   760 => x"02a9ecc0",
   761 => x"c087f2c0",
   762 => x"c002a9fb",
   763 => x"66cc87eb",
   764 => x"c703acb7",
   765 => x"0266d087",
   766 => x"537187c2",
   767 => x"c2029971",
   768 => x"fe84c187",
   769 => x"497087c3",
   770 => x"87cd0299",
   771 => x"02a9ecc0",
   772 => x"fbc087c7",
   773 => x"d5ff05a9",
   774 => x"0266d087",
   775 => x"97c087c3",
   776 => x"a9ecc07b",
   777 => x"7487c405",
   778 => x"7487c54a",
   779 => x"8a0ac04a",
   780 => x"87c24872",
   781 => x"4c264d26",
   782 => x"4f264b26",
   783 => x"87c9fd1e",
   784 => x"c04a4970",
   785 => x"c904aaf0",
   786 => x"aaf9c087",
   787 => x"c087c301",
   788 => x"c1c18af0",
   789 => x"87c904aa",
   790 => x"01aadac1",
   791 => x"f7c087c3",
   792 => x"2648728a",
   793 => x"5b5e0e4f",
   794 => x"f80e5d5c",
   795 => x"c04c7186",
   796 => x"87e0fc4d",
   797 => x"f4c04bc0",
   798 => x"49bf97c4",
   799 => x"cf04a9c0",
   800 => x"87f5fc87",
   801 => x"f4c083c1",
   802 => x"49bf97c4",
   803 => x"87f106ab",
   804 => x"97c4f4c0",
   805 => x"87cf02bf",
   806 => x"7087eefb",
   807 => x"c6029949",
   808 => x"a9ecc087",
   809 => x"c087f105",
   810 => x"87ddfb4b",
   811 => x"d8fb7e70",
   812 => x"58a6c887",
   813 => x"7087d2fb",
   814 => x"c883c14a",
   815 => x"699749a4",
   816 => x"05a96e49",
   817 => x"a4c987da",
   818 => x"49699749",
   819 => x"05a966c4",
   820 => x"a4ca87ce",
   821 => x"49699749",
   822 => x"87c405aa",
   823 => x"87d44dc1",
   824 => x"ecc0486e",
   825 => x"87c802a8",
   826 => x"fbc0486e",
   827 => x"87c405a8",
   828 => x"4dc14bc0",
   829 => x"fe029d75",
   830 => x"f3fa87ef",
   831 => x"f8487387",
   832 => x"87f0fc8e",
   833 => x"5b5e0e00",
   834 => x"f80e5d5c",
   835 => x"ff7e7186",
   836 => x"1e6e4bd4",
   837 => x"49ccdcc2",
   838 => x"c487dde9",
   839 => x"02987086",
   840 => x"c187ecc4",
   841 => x"4dbfdfde",
   842 => x"f8fc496e",
   843 => x"58a6c887",
   844 => x"c5059870",
   845 => x"48a6c487",
   846 => x"d0ff78c1",
   847 => x"c178c548",
   848 => x"66c47bd5",
   849 => x"c689c149",
   850 => x"dddec131",
   851 => x"484abf97",
   852 => x"7b70b071",
   853 => x"c448d0ff",
   854 => x"c7dcc278",
   855 => x"d049bf97",
   856 => x"87d70299",
   857 => x"d6c178c5",
   858 => x"c34ac07b",
   859 => x"82c17bff",
   860 => x"04aae0c0",
   861 => x"d0ff87f5",
   862 => x"c378c448",
   863 => x"d0ff7bff",
   864 => x"c178c548",
   865 => x"7bc17bd3",
   866 => x"b7c078c4",
   867 => x"edc206ad",
   868 => x"d4dcc287",
   869 => x"9c8d4cbf",
   870 => x"87c4c202",
   871 => x"7ed6cfc2",
   872 => x"c848a6c4",
   873 => x"c08c78c0",
   874 => x"c603acb7",
   875 => x"a4c0c887",
   876 => x"c24cc078",
   877 => x"bf97c7dc",
   878 => x"0299d049",
   879 => x"1ec087d1",
   880 => x"49ccdcc2",
   881 => x"c487e4eb",
   882 => x"4a497086",
   883 => x"c287f6c0",
   884 => x"c21ed6cf",
   885 => x"eb49ccdc",
   886 => x"86c487d1",
   887 => x"ff4a4970",
   888 => x"c5c848d0",
   889 => x"7bd4c178",
   890 => x"7bbf976e",
   891 => x"80c1486e",
   892 => x"66c47e70",
   893 => x"c888c148",
   894 => x"987058a6",
   895 => x"87e8ff05",
   896 => x"c448d0ff",
   897 => x"059a7278",
   898 => x"48c087c5",
   899 => x"c187c2c1",
   900 => x"ccdcc21e",
   901 => x"87f9e849",
   902 => x"9c7486c4",
   903 => x"87fcfd05",
   904 => x"06adb7c0",
   905 => x"dcc287d1",
   906 => x"78c048cc",
   907 => x"78c080d0",
   908 => x"dcc280f4",
   909 => x"c078bfd8",
   910 => x"fd01adb7",
   911 => x"d0ff87d3",
   912 => x"c178c548",
   913 => x"7bc07bd3",
   914 => x"48c178c4",
   915 => x"c087c2c0",
   916 => x"268ef848",
   917 => x"264c264d",
   918 => x"0e4f264b",
   919 => x"5d5c5b5e",
   920 => x"4b711e0e",
   921 => x"ab4d4cc0",
   922 => x"87e8c004",
   923 => x"1ee5f1c0",
   924 => x"c4029d75",
   925 => x"c24ac087",
   926 => x"724ac187",
   927 => x"87d0ec49",
   928 => x"7e7086c4",
   929 => x"056e84c1",
   930 => x"4c7387c2",
   931 => x"ac7385c1",
   932 => x"87d8ff06",
   933 => x"fe26486e",
   934 => x"711e87f9",
   935 => x"0566c44a",
   936 => x"497287c5",
   937 => x"2687def9",
   938 => x"5b5e0e4f",
   939 => x"1e0e5d5c",
   940 => x"de494c71",
   941 => x"f4dcc291",
   942 => x"9785714d",
   943 => x"dcc1026d",
   944 => x"e0dcc287",
   945 => x"82744abf",
   946 => x"cefe4972",
   947 => x"6e7e7087",
   948 => x"87f2c002",
   949 => x"4be8dcc2",
   950 => x"49cb4a6e",
   951 => x"87c8c7ff",
   952 => x"93cb4b74",
   953 => x"83f1dec1",
   954 => x"fcc083c4",
   955 => x"49747be1",
   956 => x"87dec1c1",
   957 => x"dec17b75",
   958 => x"49bf97de",
   959 => x"e8dcc21e",
   960 => x"87d6fe49",
   961 => x"497486c4",
   962 => x"87c6c1c1",
   963 => x"c2c149c0",
   964 => x"dcc287e5",
   965 => x"78c048c8",
   966 => x"eade49c1",
   967 => x"f2fc2687",
   968 => x"616f4c87",
   969 => x"676e6964",
   970 => x"002e2e2e",
   971 => x"5c5b5e0e",
   972 => x"4a4b710e",
   973 => x"bfe0dcc2",
   974 => x"fc497282",
   975 => x"4c7087dd",
   976 => x"87c4029c",
   977 => x"87d0e849",
   978 => x"48e0dcc2",
   979 => x"49c178c0",
   980 => x"fb87f4dd",
   981 => x"c01e87ff",
   982 => x"dac1c149",
   983 => x"1e4f2687",
   984 => x"cb494a71",
   985 => x"f1dec191",
   986 => x"1181c881",
   987 => x"ccdcc248",
   988 => x"e0dcc258",
   989 => x"c178c048",
   990 => x"87cbdd49",
   991 => x"711e4f26",
   992 => x"87d20299",
   993 => x"48c6e0c1",
   994 => x"80f750c0",
   995 => x"40dffdc0",
   996 => x"78eadec1",
   997 => x"e0c187ce",
   998 => x"dec148c2",
   999 => x"80fc78e3",
  1000 => x"78d6fdc0",
  1001 => x"5e0e4f26",
  1002 => x"0e5d5c5b",
  1003 => x"cfc286f4",
  1004 => x"4cc04dd6",
  1005 => x"c048a6c4",
  1006 => x"e0dcc278",
  1007 => x"a9c049bf",
  1008 => x"87c1c106",
  1009 => x"48d6cfc2",
  1010 => x"f8c00298",
  1011 => x"e5f1c087",
  1012 => x"0266c81e",
  1013 => x"a6c487c7",
  1014 => x"c578c048",
  1015 => x"48a6c487",
  1016 => x"66c478c1",
  1017 => x"87e8e649",
  1018 => x"4d7086c4",
  1019 => x"66c484c1",
  1020 => x"c880c148",
  1021 => x"dcc258a6",
  1022 => x"ac49bfe0",
  1023 => x"7587c603",
  1024 => x"c8ff059d",
  1025 => x"754cc087",
  1026 => x"e0c3029d",
  1027 => x"e5f1c087",
  1028 => x"0266c81e",
  1029 => x"a6cc87c7",
  1030 => x"c578c048",
  1031 => x"48a6cc87",
  1032 => x"66cc78c1",
  1033 => x"87e8e549",
  1034 => x"7e7086c4",
  1035 => x"e9c2026e",
  1036 => x"cb496e87",
  1037 => x"49699781",
  1038 => x"c10299d0",
  1039 => x"fcc087d6",
  1040 => x"49744aec",
  1041 => x"dec191cb",
  1042 => x"797281f1",
  1043 => x"ffc381c8",
  1044 => x"de497451",
  1045 => x"f4dcc291",
  1046 => x"c285714d",
  1047 => x"c17d97c1",
  1048 => x"e0c049a5",
  1049 => x"e6d7c251",
  1050 => x"d202bf97",
  1051 => x"c284c187",
  1052 => x"d7c24ba5",
  1053 => x"49db4ae6",
  1054 => x"87ecc0ff",
  1055 => x"cd87dbc1",
  1056 => x"51c049a5",
  1057 => x"a5c284c1",
  1058 => x"cb4a6e4b",
  1059 => x"d7c0ff49",
  1060 => x"87c6c187",
  1061 => x"4ae9fac0",
  1062 => x"91cb4974",
  1063 => x"81f1dec1",
  1064 => x"d7c27972",
  1065 => x"02bf97e6",
  1066 => x"497487d8",
  1067 => x"84c191de",
  1068 => x"4bf4dcc2",
  1069 => x"d7c28371",
  1070 => x"49dd4ae6",
  1071 => x"87e8fffe",
  1072 => x"4b7487d8",
  1073 => x"dcc293de",
  1074 => x"a3cb83f4",
  1075 => x"c151c049",
  1076 => x"4a6e7384",
  1077 => x"fffe49cb",
  1078 => x"66c487ce",
  1079 => x"c880c148",
  1080 => x"acc758a6",
  1081 => x"87c5c003",
  1082 => x"e0fc056e",
  1083 => x"f4487487",
  1084 => x"87dff58e",
  1085 => x"711e731e",
  1086 => x"91cb494b",
  1087 => x"81f1dec1",
  1088 => x"c14aa1c8",
  1089 => x"1248ddde",
  1090 => x"4aa1c950",
  1091 => x"48c4f4c0",
  1092 => x"81ca5012",
  1093 => x"48dedec1",
  1094 => x"dec15011",
  1095 => x"49bf97de",
  1096 => x"f549c01e",
  1097 => x"dcc287f4",
  1098 => x"78de48c8",
  1099 => x"d6d649c1",
  1100 => x"e2f42687",
  1101 => x"5b5e0e87",
  1102 => x"f40e5d5c",
  1103 => x"494d7186",
  1104 => x"dec191cb",
  1105 => x"a1c881f1",
  1106 => x"7ea1ca4a",
  1107 => x"c248a6c4",
  1108 => x"78bfd0e0",
  1109 => x"4bbf976e",
  1110 => x"734866c4",
  1111 => x"4c4b7028",
  1112 => x"a6cc4812",
  1113 => x"c19c7058",
  1114 => x"9781c984",
  1115 => x"acb74969",
  1116 => x"c087c204",
  1117 => x"bf976e4c",
  1118 => x"4966c84a",
  1119 => x"b9ff3172",
  1120 => x"749966c4",
  1121 => x"70307248",
  1122 => x"b071484a",
  1123 => x"58d4e0c2",
  1124 => x"87fee4c0",
  1125 => x"eed449c0",
  1126 => x"c0497587",
  1127 => x"f487f3f6",
  1128 => x"87eff28e",
  1129 => x"711e731e",
  1130 => x"c8fe494b",
  1131 => x"fe497387",
  1132 => x"e2f287c3",
  1133 => x"1e731e87",
  1134 => x"a3c64b71",
  1135 => x"e3c0024a",
  1136 => x"028ac187",
  1137 => x"028a87d6",
  1138 => x"8a87e8c1",
  1139 => x"87cac102",
  1140 => x"efc0028a",
  1141 => x"d9028a87",
  1142 => x"87e9c187",
  1143 => x"fef549c7",
  1144 => x"87ecc187",
  1145 => x"48c8dcc2",
  1146 => x"49c178df",
  1147 => x"c187d8d3",
  1148 => x"dcc287de",
  1149 => x"c102bfe0",
  1150 => x"c14887cb",
  1151 => x"e4dcc288",
  1152 => x"87c1c158",
  1153 => x"bfe4dcc2",
  1154 => x"87f9c002",
  1155 => x"bfe0dcc2",
  1156 => x"c280c148",
  1157 => x"c058e4dc",
  1158 => x"dcc287eb",
  1159 => x"c649bfe0",
  1160 => x"e4dcc289",
  1161 => x"a9b7c059",
  1162 => x"c287da03",
  1163 => x"c048e0dc",
  1164 => x"c287d278",
  1165 => x"02bfe4dc",
  1166 => x"dcc287cb",
  1167 => x"c648bfe0",
  1168 => x"e4dcc280",
  1169 => x"d149c058",
  1170 => x"497387fd",
  1171 => x"87c2f4c0",
  1172 => x"0e87c4f0",
  1173 => x"5d5c5b5e",
  1174 => x"86d0ff0e",
  1175 => x"c859a6dc",
  1176 => x"78c048a6",
  1177 => x"c4c180c4",
  1178 => x"80c47866",
  1179 => x"80c478c1",
  1180 => x"dcc278c1",
  1181 => x"78c148e4",
  1182 => x"bfc8dcc2",
  1183 => x"05a8de48",
  1184 => x"e1f487cb",
  1185 => x"cc497087",
  1186 => x"f9cf59a6",
  1187 => x"87c4e487",
  1188 => x"e387e6e4",
  1189 => x"4c7087f3",
  1190 => x"02acfbc0",
  1191 => x"d887fbc1",
  1192 => x"edc10566",
  1193 => x"66c0c187",
  1194 => x"6a82c44a",
  1195 => x"c11e727e",
  1196 => x"c448fbda",
  1197 => x"a1c84966",
  1198 => x"7141204a",
  1199 => x"87f905aa",
  1200 => x"4a265110",
  1201 => x"4866c0c1",
  1202 => x"78f4c3c1",
  1203 => x"81c7496a",
  1204 => x"c0c15174",
  1205 => x"81c84966",
  1206 => x"c0c151c1",
  1207 => x"81c94966",
  1208 => x"c0c151c0",
  1209 => x"81ca4966",
  1210 => x"1ec151c0",
  1211 => x"496a1ed8",
  1212 => x"d8e381c8",
  1213 => x"c186c887",
  1214 => x"c04866c4",
  1215 => x"87c701a8",
  1216 => x"c148a6c8",
  1217 => x"c187ce78",
  1218 => x"c14866c4",
  1219 => x"58a6d088",
  1220 => x"e4e287c3",
  1221 => x"48a6d087",
  1222 => x"9c7478c2",
  1223 => x"87e2cd02",
  1224 => x"c14866c8",
  1225 => x"03a866c8",
  1226 => x"dc87d7cd",
  1227 => x"78c048a6",
  1228 => x"78c080e8",
  1229 => x"7087d2e1",
  1230 => x"acd0c14c",
  1231 => x"87d7c205",
  1232 => x"e37e66c4",
  1233 => x"497087f6",
  1234 => x"e059a6c8",
  1235 => x"4c7087fb",
  1236 => x"05acecc0",
  1237 => x"c887ebc1",
  1238 => x"91cb4966",
  1239 => x"8166c0c1",
  1240 => x"6a4aa1c4",
  1241 => x"4aa1c84d",
  1242 => x"c05266c4",
  1243 => x"e079dffd",
  1244 => x"4c7087d7",
  1245 => x"87d8029c",
  1246 => x"02acfbc0",
  1247 => x"557487d2",
  1248 => x"7087c6e0",
  1249 => x"c7029c4c",
  1250 => x"acfbc087",
  1251 => x"87eeff05",
  1252 => x"c255e0c0",
  1253 => x"97c055c1",
  1254 => x"4966d87d",
  1255 => x"db05a96e",
  1256 => x"4866c887",
  1257 => x"04a866cc",
  1258 => x"66c887ca",
  1259 => x"cc80c148",
  1260 => x"87c858a6",
  1261 => x"c14866cc",
  1262 => x"58a6d088",
  1263 => x"87c9dfff",
  1264 => x"d0c14c70",
  1265 => x"87c805ac",
  1266 => x"c14866d4",
  1267 => x"58a6d880",
  1268 => x"02acd0c1",
  1269 => x"c087e9fd",
  1270 => x"d848a6e0",
  1271 => x"66c47866",
  1272 => x"66e0c048",
  1273 => x"ebc905a8",
  1274 => x"a6e4c087",
  1275 => x"7478c048",
  1276 => x"88fbc048",
  1277 => x"026e7e70",
  1278 => x"6e87eec9",
  1279 => x"7088cb48",
  1280 => x"c1026e7e",
  1281 => x"486e87cd",
  1282 => x"7e7088c9",
  1283 => x"c1c4026e",
  1284 => x"c4486e87",
  1285 => x"6e7e7088",
  1286 => x"6e87ce02",
  1287 => x"7088c148",
  1288 => x"c3026e7e",
  1289 => x"e2c887ec",
  1290 => x"48a6dc87",
  1291 => x"ff78f0c0",
  1292 => x"7087d6dd",
  1293 => x"acecc04c",
  1294 => x"87c4c002",
  1295 => x"5ca6e0c0",
  1296 => x"02acecc0",
  1297 => x"dcff87cd",
  1298 => x"4c7087ff",
  1299 => x"05acecc0",
  1300 => x"c087f3ff",
  1301 => x"c002acec",
  1302 => x"dcff87c4",
  1303 => x"1ec087eb",
  1304 => x"66d01eca",
  1305 => x"c191cb49",
  1306 => x"714866c8",
  1307 => x"58a6cc80",
  1308 => x"c44866c8",
  1309 => x"58a6d080",
  1310 => x"49bf66cc",
  1311 => x"87cdddff",
  1312 => x"1ede1ec1",
  1313 => x"49bf66d4",
  1314 => x"87c1ddff",
  1315 => x"497086d0",
  1316 => x"c08909c0",
  1317 => x"c059a6ec",
  1318 => x"c04866e8",
  1319 => x"eec006a8",
  1320 => x"66e8c087",
  1321 => x"03a8dd48",
  1322 => x"c487e4c0",
  1323 => x"c049bf66",
  1324 => x"c08166e8",
  1325 => x"e8c051e0",
  1326 => x"81c14966",
  1327 => x"81bf66c4",
  1328 => x"c051c1c2",
  1329 => x"c24966e8",
  1330 => x"bf66c481",
  1331 => x"6e51c081",
  1332 => x"f4c3c148",
  1333 => x"c8496e78",
  1334 => x"5166d081",
  1335 => x"81c9496e",
  1336 => x"6e5166d4",
  1337 => x"dc81ca49",
  1338 => x"66d05166",
  1339 => x"d480c148",
  1340 => x"66c858a6",
  1341 => x"a866cc48",
  1342 => x"87cbc004",
  1343 => x"c14866c8",
  1344 => x"58a6cc80",
  1345 => x"cc87e2c5",
  1346 => x"88c14866",
  1347 => x"c558a6d0",
  1348 => x"dcff87d7",
  1349 => x"497087e6",
  1350 => x"59a6ecc0",
  1351 => x"87dcdcff",
  1352 => x"e0c04970",
  1353 => x"66dc59a6",
  1354 => x"a8ecc048",
  1355 => x"87cac005",
  1356 => x"c048a6dc",
  1357 => x"c07866e8",
  1358 => x"d9ff87c4",
  1359 => x"66c887cb",
  1360 => x"c191cb49",
  1361 => x"714866c0",
  1362 => x"6e7e7080",
  1363 => x"6e82c84a",
  1364 => x"c081ca49",
  1365 => x"dc5166e8",
  1366 => x"81c14966",
  1367 => x"8966e8c0",
  1368 => x"307148c1",
  1369 => x"89c14970",
  1370 => x"c27a9771",
  1371 => x"49bfd0e0",
  1372 => x"2966e8c0",
  1373 => x"484a6a97",
  1374 => x"f0c09871",
  1375 => x"496e58a6",
  1376 => x"4d6981c4",
  1377 => x"4866e0c0",
  1378 => x"02a866c4",
  1379 => x"c487c8c0",
  1380 => x"78c048a6",
  1381 => x"c487c5c0",
  1382 => x"78c148a6",
  1383 => x"c01e66c4",
  1384 => x"49751ee0",
  1385 => x"87e5d8ff",
  1386 => x"4c7086c8",
  1387 => x"06acb7c0",
  1388 => x"7487d4c1",
  1389 => x"49e0c085",
  1390 => x"4b758974",
  1391 => x"4ac4dbc1",
  1392 => x"e3ebfe71",
  1393 => x"c085c287",
  1394 => x"c14866e4",
  1395 => x"a6e8c080",
  1396 => x"66ecc058",
  1397 => x"7081c149",
  1398 => x"c8c002a9",
  1399 => x"48a6c487",
  1400 => x"c5c078c0",
  1401 => x"48a6c487",
  1402 => x"66c478c1",
  1403 => x"49a4c21e",
  1404 => x"7148e0c0",
  1405 => x"1e497088",
  1406 => x"d7ff4975",
  1407 => x"86c887cf",
  1408 => x"01a8b7c0",
  1409 => x"c087c0ff",
  1410 => x"c00266e4",
  1411 => x"496e87d1",
  1412 => x"e4c081c9",
  1413 => x"486e5166",
  1414 => x"78f5c4c1",
  1415 => x"6e87ccc0",
  1416 => x"c281c949",
  1417 => x"c1486e51",
  1418 => x"c878e4c6",
  1419 => x"66cc4866",
  1420 => x"cbc004a8",
  1421 => x"4866c887",
  1422 => x"a6cc80c1",
  1423 => x"87e9c058",
  1424 => x"c14866cc",
  1425 => x"58a6d088",
  1426 => x"ff87dec0",
  1427 => x"7087ead5",
  1428 => x"87d5c04c",
  1429 => x"05acc6c1",
  1430 => x"d087c8c0",
  1431 => x"80c14866",
  1432 => x"ff58a6d4",
  1433 => x"7087d2d5",
  1434 => x"4866d44c",
  1435 => x"a6d880c1",
  1436 => x"029c7458",
  1437 => x"c887cbc0",
  1438 => x"c8c14866",
  1439 => x"f204a866",
  1440 => x"d4ff87e9",
  1441 => x"66c887ea",
  1442 => x"03a8c748",
  1443 => x"c287e5c0",
  1444 => x"c048e4dc",
  1445 => x"4966c878",
  1446 => x"c0c191cb",
  1447 => x"a1c48166",
  1448 => x"c04a6a4a",
  1449 => x"66c87952",
  1450 => x"cc80c148",
  1451 => x"a8c758a6",
  1452 => x"87dbff04",
  1453 => x"ff8ed0ff",
  1454 => x"4c87d8de",
  1455 => x"2064616f",
  1456 => x"00202e2a",
  1457 => x"1e00203a",
  1458 => x"4b711e73",
  1459 => x"87c6029b",
  1460 => x"48e0dcc2",
  1461 => x"1ec778c0",
  1462 => x"bfe0dcc2",
  1463 => x"dec11e49",
  1464 => x"dcc21ef1",
  1465 => x"ed49bfc8",
  1466 => x"86cc87e9",
  1467 => x"bfc8dcc2",
  1468 => x"87cae249",
  1469 => x"c8029b73",
  1470 => x"f1dec187",
  1471 => x"e3e2c049",
  1472 => x"d2ddff87",
  1473 => x"dec11e87",
  1474 => x"50c048dd",
  1475 => x"bfd4e0c1",
  1476 => x"f0d7ff49",
  1477 => x"2648c087",
  1478 => x"dec71e4f",
  1479 => x"fe49c187",
  1480 => x"eefe87e5",
  1481 => x"987087c3",
  1482 => x"fe87cd02",
  1483 => x"7087dcf5",
  1484 => x"87c40298",
  1485 => x"87c24ac1",
  1486 => x"9a724ac0",
  1487 => x"c087ce05",
  1488 => x"f4ddc11e",
  1489 => x"e0efc049",
  1490 => x"fe86c487",
  1491 => x"e0dcc287",
  1492 => x"c278c048",
  1493 => x"c048c8dc",
  1494 => x"ddc11e78",
  1495 => x"efc049ff",
  1496 => x"1ec087c7",
  1497 => x"7087defe",
  1498 => x"fceec049",
  1499 => x"87cac387",
  1500 => x"4f268ef8",
  1501 => x"66204453",
  1502 => x"656c6961",
  1503 => x"42002e64",
  1504 => x"69746f6f",
  1505 => x"2e2e676e",
  1506 => x"c01e002e",
  1507 => x"fa87d2e2",
  1508 => x"1e4f2687",
  1509 => x"f187c2fe",
  1510 => x"2648c087",
  1511 => x"0100004f",
  1512 => x"80000000",
  1513 => x"69784520",
  1514 => x"20800074",
  1515 => x"6b636142",
  1516 => x"000ea900",
  1517 => x"00273400",
  1518 => x"00000000",
  1519 => x"00000ea9",
  1520 => x"00002752",
  1521 => x"a9000000",
  1522 => x"7000000e",
  1523 => x"00000027",
  1524 => x"0ea90000",
  1525 => x"278e0000",
  1526 => x"00000000",
  1527 => x"000ea900",
  1528 => x"0027ac00",
  1529 => x"00000000",
  1530 => x"00000ea9",
  1531 => x"000027ca",
  1532 => x"a9000000",
  1533 => x"e800000e",
  1534 => x"00000027",
  1535 => x"0f5f0000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"0011b500",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00001818",
  1542 => x"544f4f42",
  1543 => x"20202020",
  1544 => x"004d4f52",
  1545 => x"48f0fe1e",
  1546 => x"09cd78c0",
  1547 => x"4f260979",
  1548 => x"f0fe1e1e",
  1549 => x"26487ebf",
  1550 => x"fe1e4f26",
  1551 => x"78c148f0",
  1552 => x"fe1e4f26",
  1553 => x"78c048f0",
  1554 => x"711e4f26",
  1555 => x"5252c04a",
  1556 => x"5e0e4f26",
  1557 => x"0e5d5c5b",
  1558 => x"4d7186f4",
  1559 => x"c17e6d97",
  1560 => x"6c974ca5",
  1561 => x"58a6c848",
  1562 => x"66c4486e",
  1563 => x"87c505a8",
  1564 => x"e6c048ff",
  1565 => x"87caff87",
  1566 => x"9749a5c2",
  1567 => x"a3714b6c",
  1568 => x"4b6b974b",
  1569 => x"6e7e6c97",
  1570 => x"c880c148",
  1571 => x"98c758a6",
  1572 => x"7058a6cc",
  1573 => x"e1fe7c97",
  1574 => x"f4487387",
  1575 => x"264d268e",
  1576 => x"264b264c",
  1577 => x"5b5e0e4f",
  1578 => x"86f40e5c",
  1579 => x"66d84c71",
  1580 => x"9affc34a",
  1581 => x"974ba4c2",
  1582 => x"a173496c",
  1583 => x"97517249",
  1584 => x"486e7e6c",
  1585 => x"a6c880c1",
  1586 => x"cc98c758",
  1587 => x"547058a6",
  1588 => x"caff8ef4",
  1589 => x"fd1e1e87",
  1590 => x"bfe087e8",
  1591 => x"e0c0494a",
  1592 => x"cb0299c0",
  1593 => x"c21e7287",
  1594 => x"fe49c6e0",
  1595 => x"86c487f7",
  1596 => x"7087fdfc",
  1597 => x"87c2fd7e",
  1598 => x"1e4f2626",
  1599 => x"49c6e0c2",
  1600 => x"c187c7fd",
  1601 => x"fc49d5e3",
  1602 => x"eec387da",
  1603 => x"0e4f2687",
  1604 => x"5d5c5b5e",
  1605 => x"c24d710e",
  1606 => x"fc49c6e0",
  1607 => x"4b7087f4",
  1608 => x"04abb7c0",
  1609 => x"c387c2c3",
  1610 => x"c905abf0",
  1611 => x"f3e7c187",
  1612 => x"c278c148",
  1613 => x"e0c387e3",
  1614 => x"87c905ab",
  1615 => x"48f7e7c1",
  1616 => x"d4c278c1",
  1617 => x"f7e7c187",
  1618 => x"87c602bf",
  1619 => x"4ca3c0c2",
  1620 => x"4c7387c2",
  1621 => x"bff3e7c1",
  1622 => x"87e0c002",
  1623 => x"b7c44974",
  1624 => x"e9c19129",
  1625 => x"4a7481ca",
  1626 => x"92c29acf",
  1627 => x"307248c1",
  1628 => x"baff4a70",
  1629 => x"98694872",
  1630 => x"87db7970",
  1631 => x"b7c44974",
  1632 => x"e9c19129",
  1633 => x"4a7481ca",
  1634 => x"92c29acf",
  1635 => x"307248c3",
  1636 => x"69484a70",
  1637 => x"757970b0",
  1638 => x"f0c0059d",
  1639 => x"48d0ff87",
  1640 => x"ff78e1c8",
  1641 => x"78c548d4",
  1642 => x"bff7e7c1",
  1643 => x"c387c302",
  1644 => x"e7c178e0",
  1645 => x"c602bff3",
  1646 => x"48d4ff87",
  1647 => x"ff78f0c3",
  1648 => x"787348d4",
  1649 => x"c848d0ff",
  1650 => x"e0c078e1",
  1651 => x"f7e7c178",
  1652 => x"c178c048",
  1653 => x"c048f3e7",
  1654 => x"c6e0c278",
  1655 => x"87f2f949",
  1656 => x"b7c04b70",
  1657 => x"fefc03ab",
  1658 => x"2648c087",
  1659 => x"264c264d",
  1660 => x"004f264b",
  1661 => x"00000000",
  1662 => x"1e000000",
  1663 => x"49724ac0",
  1664 => x"e9c191c4",
  1665 => x"79c081ca",
  1666 => x"b7d082c1",
  1667 => x"87ee04aa",
  1668 => x"5e0e4f26",
  1669 => x"0e5d5c5b",
  1670 => x"e5f84d71",
  1671 => x"c44a7587",
  1672 => x"c1922ab7",
  1673 => x"7582cae9",
  1674 => x"c29ccf4c",
  1675 => x"4b496a94",
  1676 => x"9bc32b74",
  1677 => x"307448c2",
  1678 => x"bcff4c70",
  1679 => x"98714874",
  1680 => x"f5f77a70",
  1681 => x"fe487387",
  1682 => x"000087e1",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"ff1e0000",
  1699 => x"e1c848d0",
  1700 => x"ff487178",
  1701 => x"c47808d4",
  1702 => x"d4ff4866",
  1703 => x"4f267808",
  1704 => x"c44a711e",
  1705 => x"721e4966",
  1706 => x"87deff49",
  1707 => x"c048d0ff",
  1708 => x"262678e0",
  1709 => x"1e731e4f",
  1710 => x"66c84b71",
  1711 => x"4a731e49",
  1712 => x"49a2e0c1",
  1713 => x"2687d9ff",
  1714 => x"4d2687c4",
  1715 => x"4b264c26",
  1716 => x"ff1e4f26",
  1717 => x"ffc34ad4",
  1718 => x"48d0ff7a",
  1719 => x"de78e1c0",
  1720 => x"d0e0c27a",
  1721 => x"48497abf",
  1722 => x"7a7028c8",
  1723 => x"28d04871",
  1724 => x"48717a70",
  1725 => x"7a7028d8",
  1726 => x"c048d0ff",
  1727 => x"4f2678e0",
  1728 => x"48d0ff1e",
  1729 => x"7178c9c8",
  1730 => x"08d4ff48",
  1731 => x"1e4f2678",
  1732 => x"eb494a71",
  1733 => x"48d0ff87",
  1734 => x"4f2678c8",
  1735 => x"711e731e",
  1736 => x"e0e0c24b",
  1737 => x"87c302bf",
  1738 => x"ff87ebc2",
  1739 => x"c9c848d0",
  1740 => x"c0497378",
  1741 => x"d4ffb1e0",
  1742 => x"c2787148",
  1743 => x"c048d4e0",
  1744 => x"0266c878",
  1745 => x"ffc387c5",
  1746 => x"c087c249",
  1747 => x"dce0c249",
  1748 => x"0266cc59",
  1749 => x"d5c587c6",
  1750 => x"87c44ad5",
  1751 => x"4affffcf",
  1752 => x"5ae0e0c2",
  1753 => x"48e0e0c2",
  1754 => x"87c478c1",
  1755 => x"4c264d26",
  1756 => x"4f264b26",
  1757 => x"5c5b5e0e",
  1758 => x"4a710e5d",
  1759 => x"bfdce0c2",
  1760 => x"029a724c",
  1761 => x"c84987cb",
  1762 => x"d2ecc191",
  1763 => x"c483714b",
  1764 => x"d2f0c187",
  1765 => x"134dc04b",
  1766 => x"c2997449",
  1767 => x"b9bfd8e0",
  1768 => x"7148d4ff",
  1769 => x"2cb7c178",
  1770 => x"adb7c885",
  1771 => x"c287e804",
  1772 => x"48bfd4e0",
  1773 => x"e0c280c8",
  1774 => x"effe58d8",
  1775 => x"1e731e87",
  1776 => x"4a134b71",
  1777 => x"87cb029a",
  1778 => x"e7fe4972",
  1779 => x"9a4a1387",
  1780 => x"fe87f505",
  1781 => x"c21e87da",
  1782 => x"49bfd4e0",
  1783 => x"48d4e0c2",
  1784 => x"c478a1c1",
  1785 => x"03a9b7c0",
  1786 => x"d4ff87db",
  1787 => x"d8e0c248",
  1788 => x"e0c278bf",
  1789 => x"c249bfd4",
  1790 => x"c148d4e0",
  1791 => x"c0c478a1",
  1792 => x"e504a9b7",
  1793 => x"48d0ff87",
  1794 => x"e0c278c8",
  1795 => x"78c048e0",
  1796 => x"00004f26",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"005f5f00",
  1800 => x"03000000",
  1801 => x"03030003",
  1802 => x"7f140000",
  1803 => x"7f7f147f",
  1804 => x"24000014",
  1805 => x"3a6b6b2e",
  1806 => x"6a4c0012",
  1807 => x"566c1836",
  1808 => x"7e300032",
  1809 => x"3a77594f",
  1810 => x"00004068",
  1811 => x"00030704",
  1812 => x"00000000",
  1813 => x"41633e1c",
  1814 => x"00000000",
  1815 => x"1c3e6341",
  1816 => x"2a080000",
  1817 => x"3e1c1c3e",
  1818 => x"0800082a",
  1819 => x"083e3e08",
  1820 => x"00000008",
  1821 => x"0060e080",
  1822 => x"08000000",
  1823 => x"08080808",
  1824 => x"00000008",
  1825 => x"00606000",
  1826 => x"60400000",
  1827 => x"060c1830",
  1828 => x"3e000103",
  1829 => x"7f4d597f",
  1830 => x"0400003e",
  1831 => x"007f7f06",
  1832 => x"42000000",
  1833 => x"4f597163",
  1834 => x"22000046",
  1835 => x"7f494963",
  1836 => x"1c180036",
  1837 => x"7f7f1316",
  1838 => x"27000010",
  1839 => x"7d454567",
  1840 => x"3c000039",
  1841 => x"79494b7e",
  1842 => x"01000030",
  1843 => x"0f797101",
  1844 => x"36000007",
  1845 => x"7f49497f",
  1846 => x"06000036",
  1847 => x"3f69494f",
  1848 => x"0000001e",
  1849 => x"00666600",
  1850 => x"00000000",
  1851 => x"0066e680",
  1852 => x"08000000",
  1853 => x"22141408",
  1854 => x"14000022",
  1855 => x"14141414",
  1856 => x"22000014",
  1857 => x"08141422",
  1858 => x"02000008",
  1859 => x"0f595103",
  1860 => x"7f3e0006",
  1861 => x"1f555d41",
  1862 => x"7e00001e",
  1863 => x"7f09097f",
  1864 => x"7f00007e",
  1865 => x"7f49497f",
  1866 => x"1c000036",
  1867 => x"4141633e",
  1868 => x"7f000041",
  1869 => x"3e63417f",
  1870 => x"7f00001c",
  1871 => x"4149497f",
  1872 => x"7f000041",
  1873 => x"0109097f",
  1874 => x"3e000001",
  1875 => x"7b49417f",
  1876 => x"7f00007a",
  1877 => x"7f08087f",
  1878 => x"0000007f",
  1879 => x"417f7f41",
  1880 => x"20000000",
  1881 => x"7f404060",
  1882 => x"7f7f003f",
  1883 => x"63361c08",
  1884 => x"7f000041",
  1885 => x"4040407f",
  1886 => x"7f7f0040",
  1887 => x"7f060c06",
  1888 => x"7f7f007f",
  1889 => x"7f180c06",
  1890 => x"3e00007f",
  1891 => x"7f41417f",
  1892 => x"7f00003e",
  1893 => x"0f09097f",
  1894 => x"7f3e0006",
  1895 => x"7e7f6141",
  1896 => x"7f000040",
  1897 => x"7f19097f",
  1898 => x"26000066",
  1899 => x"7b594d6f",
  1900 => x"01000032",
  1901 => x"017f7f01",
  1902 => x"3f000001",
  1903 => x"7f40407f",
  1904 => x"0f00003f",
  1905 => x"3f70703f",
  1906 => x"7f7f000f",
  1907 => x"7f301830",
  1908 => x"6341007f",
  1909 => x"361c1c36",
  1910 => x"03014163",
  1911 => x"067c7c06",
  1912 => x"71610103",
  1913 => x"43474d59",
  1914 => x"00000041",
  1915 => x"41417f7f",
  1916 => x"03010000",
  1917 => x"30180c06",
  1918 => x"00004060",
  1919 => x"7f7f4141",
  1920 => x"0c080000",
  1921 => x"0c060306",
  1922 => x"80800008",
  1923 => x"80808080",
  1924 => x"00000080",
  1925 => x"04070300",
  1926 => x"20000000",
  1927 => x"7c545474",
  1928 => x"7f000078",
  1929 => x"7c44447f",
  1930 => x"38000038",
  1931 => x"4444447c",
  1932 => x"38000000",
  1933 => x"7f44447c",
  1934 => x"3800007f",
  1935 => x"5c54547c",
  1936 => x"04000018",
  1937 => x"05057f7e",
  1938 => x"18000000",
  1939 => x"fca4a4bc",
  1940 => x"7f00007c",
  1941 => x"7c04047f",
  1942 => x"00000078",
  1943 => x"407d3d00",
  1944 => x"80000000",
  1945 => x"7dfd8080",
  1946 => x"7f000000",
  1947 => x"6c38107f",
  1948 => x"00000044",
  1949 => x"407f3f00",
  1950 => x"7c7c0000",
  1951 => x"7c0c180c",
  1952 => x"7c000078",
  1953 => x"7c04047c",
  1954 => x"38000078",
  1955 => x"7c44447c",
  1956 => x"fc000038",
  1957 => x"3c2424fc",
  1958 => x"18000018",
  1959 => x"fc24243c",
  1960 => x"7c0000fc",
  1961 => x"0c04047c",
  1962 => x"48000008",
  1963 => x"7454545c",
  1964 => x"04000020",
  1965 => x"44447f3f",
  1966 => x"3c000000",
  1967 => x"7c40407c",
  1968 => x"1c00007c",
  1969 => x"3c60603c",
  1970 => x"7c3c001c",
  1971 => x"7c603060",
  1972 => x"6c44003c",
  1973 => x"6c381038",
  1974 => x"1c000044",
  1975 => x"3c60e0bc",
  1976 => x"4400001c",
  1977 => x"4c5c7464",
  1978 => x"08000044",
  1979 => x"41773e08",
  1980 => x"00000041",
  1981 => x"007f7f00",
  1982 => x"41000000",
  1983 => x"083e7741",
  1984 => x"01020008",
  1985 => x"02020301",
  1986 => x"7f7f0001",
  1987 => x"7f7f7f7f",
  1988 => x"0808007f",
  1989 => x"3e3e1c1c",
  1990 => x"7f7f7f7f",
  1991 => x"1c1c3e3e",
  1992 => x"10000808",
  1993 => x"187c7c18",
  1994 => x"10000010",
  1995 => x"307c7c30",
  1996 => x"30100010",
  1997 => x"1e786060",
  1998 => x"66420006",
  1999 => x"663c183c",
  2000 => x"38780042",
  2001 => x"6cc6c26a",
  2002 => x"00600038",
  2003 => x"00006000",
  2004 => x"5e0e0060",
  2005 => x"0e5d5c5b",
  2006 => x"c24c711e",
  2007 => x"4dbfe5e0",
  2008 => x"1ec04bc0",
  2009 => x"c702ab74",
  2010 => x"48a6c487",
  2011 => x"87c578c0",
  2012 => x"c148a6c4",
  2013 => x"1e66c478",
  2014 => x"dfee4973",
  2015 => x"c086c887",
  2016 => x"efef49e0",
  2017 => x"4aa5c487",
  2018 => x"f0f0496a",
  2019 => x"87c6f187",
  2020 => x"83c185cb",
  2021 => x"04abb7c8",
  2022 => x"2687c7ff",
  2023 => x"4c264d26",
  2024 => x"4f264b26",
  2025 => x"c24a711e",
  2026 => x"c25ae9e0",
  2027 => x"c748e9e0",
  2028 => x"ddfe4978",
  2029 => x"1e4f2687",
  2030 => x"4a711e73",
  2031 => x"03aab7c0",
  2032 => x"cec287d3",
  2033 => x"c405bfc2",
  2034 => x"c24bc187",
  2035 => x"c24bc087",
  2036 => x"c45bc6ce",
  2037 => x"c6cec287",
  2038 => x"c2cec25a",
  2039 => x"9ac14abf",
  2040 => x"49a2c0c1",
  2041 => x"fc87e8ec",
  2042 => x"c2cec248",
  2043 => x"effe78bf",
  2044 => x"4a711e87",
  2045 => x"721e66c4",
  2046 => x"87f9ea49",
  2047 => x"1e4f2626",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
