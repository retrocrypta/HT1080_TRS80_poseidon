
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"e0",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f0",x"e0",x"c2"),
    14 => (x"48",x"f0",x"ce",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c8",x"dd"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d6",x"02",x"99",x"71"),
    50 => (x"48",x"d4",x"ff",x"87"),
    51 => (x"68",x"78",x"ff",x"c3"),
    52 => (x"49",x"66",x"c4",x"52"),
    53 => (x"c8",x"88",x"c1",x"48"),
    54 => (x"99",x"71",x"58",x"a6"),
    55 => (x"26",x"87",x"ea",x"05"),
    56 => (x"1e",x"73",x"1e",x"4f"),
    57 => (x"c3",x"4b",x"d4",x"ff"),
    58 => (x"4a",x"6b",x"7b",x"ff"),
    59 => (x"6b",x"7b",x"ff",x"c3"),
    60 => (x"72",x"32",x"c8",x"49"),
    61 => (x"7b",x"ff",x"c3",x"b1"),
    62 => (x"31",x"c8",x"4a",x"6b"),
    63 => (x"ff",x"c3",x"b2",x"71"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"71",x"b1",x"72",x"32"),
    66 => (x"26",x"87",x"c4",x"48"),
    67 => (x"26",x"4c",x"26",x"4d"),
    68 => (x"0e",x"4f",x"26",x"4b"),
    69 => (x"5d",x"5c",x"5b",x"5e"),
    70 => (x"ff",x"4a",x"71",x"0e"),
    71 => (x"49",x"72",x"4c",x"d4"),
    72 => (x"71",x"99",x"ff",x"c3"),
    73 => (x"f0",x"ce",x"c2",x"7c"),
    74 => (x"87",x"c8",x"05",x"bf"),
    75 => (x"c9",x"48",x"66",x"d0"),
    76 => (x"58",x"a6",x"d4",x"30"),
    77 => (x"d8",x"49",x"66",x"d0"),
    78 => (x"99",x"ff",x"c3",x"29"),
    79 => (x"66",x"d0",x"7c",x"71"),
    80 => (x"c3",x"29",x"d0",x"49"),
    81 => (x"7c",x"71",x"99",x"ff"),
    82 => (x"c8",x"49",x"66",x"d0"),
    83 => (x"99",x"ff",x"c3",x"29"),
    84 => (x"66",x"d0",x"7c",x"71"),
    85 => (x"99",x"ff",x"c3",x"49"),
    86 => (x"49",x"72",x"7c",x"71"),
    87 => (x"ff",x"c3",x"29",x"d0"),
    88 => (x"6c",x"7c",x"71",x"99"),
    89 => (x"ff",x"f0",x"c9",x"4b"),
    90 => (x"ab",x"ff",x"c3",x"4d"),
    91 => (x"c3",x"87",x"d0",x"05"),
    92 => (x"4b",x"6c",x"7c",x"ff"),
    93 => (x"c6",x"02",x"8d",x"c1"),
    94 => (x"ab",x"ff",x"c3",x"87"),
    95 => (x"73",x"87",x"f0",x"02"),
    96 => (x"87",x"c7",x"fe",x"48"),
    97 => (x"ff",x"49",x"c0",x"1e"),
    98 => (x"ff",x"c3",x"48",x"d4"),
    99 => (x"c3",x"81",x"c1",x"78"),
   100 => (x"04",x"a9",x"b7",x"c8"),
   101 => (x"4f",x"26",x"87",x"f1"),
   102 => (x"e7",x"1e",x"73",x"1e"),
   103 => (x"df",x"f8",x"c4",x"87"),
   104 => (x"c0",x"1e",x"c0",x"4b"),
   105 => (x"f7",x"c1",x"f0",x"ff"),
   106 => (x"87",x"e7",x"fd",x"49"),
   107 => (x"a8",x"c1",x"86",x"c4"),
   108 => (x"87",x"ea",x"c0",x"05"),
   109 => (x"c3",x"48",x"d4",x"ff"),
   110 => (x"c0",x"c1",x"78",x"ff"),
   111 => (x"c0",x"c0",x"c0",x"c0"),
   112 => (x"f0",x"e1",x"c0",x"1e"),
   113 => (x"fd",x"49",x"e9",x"c1"),
   114 => (x"86",x"c4",x"87",x"c9"),
   115 => (x"ca",x"05",x"98",x"70"),
   116 => (x"48",x"d4",x"ff",x"87"),
   117 => (x"c1",x"78",x"ff",x"c3"),
   118 => (x"fe",x"87",x"cb",x"48"),
   119 => (x"8b",x"c1",x"87",x"e6"),
   120 => (x"87",x"fd",x"fe",x"05"),
   121 => (x"e6",x"fc",x"48",x"c0"),
   122 => (x"1e",x"73",x"1e",x"87"),
   123 => (x"c3",x"48",x"d4",x"ff"),
   124 => (x"4b",x"d3",x"78",x"ff"),
   125 => (x"ff",x"c0",x"1e",x"c0"),
   126 => (x"49",x"c1",x"c1",x"f0"),
   127 => (x"c4",x"87",x"d4",x"fc"),
   128 => (x"05",x"98",x"70",x"86"),
   129 => (x"d4",x"ff",x"87",x"ca"),
   130 => (x"78",x"ff",x"c3",x"48"),
   131 => (x"87",x"cb",x"48",x"c1"),
   132 => (x"c1",x"87",x"f1",x"fd"),
   133 => (x"db",x"ff",x"05",x"8b"),
   134 => (x"fb",x"48",x"c0",x"87"),
   135 => (x"5e",x"0e",x"87",x"f1"),
   136 => (x"ff",x"0e",x"5c",x"5b"),
   137 => (x"db",x"fd",x"4c",x"d4"),
   138 => (x"1e",x"ea",x"c6",x"87"),
   139 => (x"c1",x"f0",x"e1",x"c0"),
   140 => (x"de",x"fb",x"49",x"c8"),
   141 => (x"c1",x"86",x"c4",x"87"),
   142 => (x"87",x"c8",x"02",x"a8"),
   143 => (x"c0",x"87",x"ea",x"fe"),
   144 => (x"87",x"e2",x"c1",x"48"),
   145 => (x"70",x"87",x"da",x"fa"),
   146 => (x"ff",x"ff",x"cf",x"49"),
   147 => (x"a9",x"ea",x"c6",x"99"),
   148 => (x"fe",x"87",x"c8",x"02"),
   149 => (x"48",x"c0",x"87",x"d3"),
   150 => (x"c3",x"87",x"cb",x"c1"),
   151 => (x"f1",x"c0",x"7c",x"ff"),
   152 => (x"87",x"f4",x"fc",x"4b"),
   153 => (x"c0",x"02",x"98",x"70"),
   154 => (x"1e",x"c0",x"87",x"eb"),
   155 => (x"c1",x"f0",x"ff",x"c0"),
   156 => (x"de",x"fa",x"49",x"fa"),
   157 => (x"70",x"86",x"c4",x"87"),
   158 => (x"87",x"d9",x"05",x"98"),
   159 => (x"6c",x"7c",x"ff",x"c3"),
   160 => (x"7c",x"ff",x"c3",x"49"),
   161 => (x"c1",x"7c",x"7c",x"7c"),
   162 => (x"c4",x"02",x"99",x"c0"),
   163 => (x"d5",x"48",x"c1",x"87"),
   164 => (x"d1",x"48",x"c0",x"87"),
   165 => (x"05",x"ab",x"c2",x"87"),
   166 => (x"48",x"c0",x"87",x"c4"),
   167 => (x"8b",x"c1",x"87",x"c8"),
   168 => (x"87",x"fd",x"fe",x"05"),
   169 => (x"e4",x"f9",x"48",x"c0"),
   170 => (x"1e",x"73",x"1e",x"87"),
   171 => (x"48",x"f0",x"ce",x"c2"),
   172 => (x"4b",x"c7",x"78",x"c1"),
   173 => (x"c2",x"48",x"d0",x"ff"),
   174 => (x"87",x"c8",x"fb",x"78"),
   175 => (x"c3",x"48",x"d0",x"ff"),
   176 => (x"c0",x"1e",x"c0",x"78"),
   177 => (x"c0",x"c1",x"d0",x"e5"),
   178 => (x"87",x"c7",x"f9",x"49"),
   179 => (x"a8",x"c1",x"86",x"c4"),
   180 => (x"4b",x"87",x"c1",x"05"),
   181 => (x"c5",x"05",x"ab",x"c2"),
   182 => (x"c0",x"48",x"c0",x"87"),
   183 => (x"8b",x"c1",x"87",x"f9"),
   184 => (x"87",x"d0",x"ff",x"05"),
   185 => (x"c2",x"87",x"f7",x"fc"),
   186 => (x"70",x"58",x"f4",x"ce"),
   187 => (x"87",x"cd",x"05",x"98"),
   188 => (x"ff",x"c0",x"1e",x"c1"),
   189 => (x"49",x"d0",x"c1",x"f0"),
   190 => (x"c4",x"87",x"d8",x"f8"),
   191 => (x"48",x"d4",x"ff",x"86"),
   192 => (x"c2",x"78",x"ff",x"c3"),
   193 => (x"ce",x"c2",x"87",x"fc"),
   194 => (x"d0",x"ff",x"58",x"f8"),
   195 => (x"ff",x"78",x"c2",x"48"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"f7",x"48",x"c1",x"78"),
   198 => (x"5e",x"0e",x"87",x"f5"),
   199 => (x"0e",x"5d",x"5c",x"5b"),
   200 => (x"4c",x"c0",x"4b",x"71"),
   201 => (x"df",x"cd",x"ee",x"c5"),
   202 => (x"48",x"d4",x"ff",x"4a"),
   203 => (x"68",x"78",x"ff",x"c3"),
   204 => (x"a9",x"fe",x"c3",x"49"),
   205 => (x"87",x"fd",x"c0",x"05"),
   206 => (x"9b",x"73",x"4d",x"70"),
   207 => (x"d0",x"87",x"cc",x"02"),
   208 => (x"49",x"73",x"1e",x"66"),
   209 => (x"c4",x"87",x"f1",x"f5"),
   210 => (x"ff",x"87",x"d6",x"86"),
   211 => (x"d1",x"c4",x"48",x"d0"),
   212 => (x"7d",x"ff",x"c3",x"78"),
   213 => (x"c1",x"48",x"66",x"d0"),
   214 => (x"58",x"a6",x"d4",x"88"),
   215 => (x"f0",x"05",x"98",x"70"),
   216 => (x"48",x"d4",x"ff",x"87"),
   217 => (x"78",x"78",x"ff",x"c3"),
   218 => (x"c5",x"05",x"9b",x"73"),
   219 => (x"48",x"d0",x"ff",x"87"),
   220 => (x"4a",x"c1",x"78",x"d0"),
   221 => (x"05",x"8a",x"c1",x"4c"),
   222 => (x"74",x"87",x"ee",x"fe"),
   223 => (x"87",x"cb",x"f6",x"48"),
   224 => (x"71",x"1e",x"73",x"1e"),
   225 => (x"ff",x"4b",x"c0",x"4a"),
   226 => (x"ff",x"c3",x"48",x"d4"),
   227 => (x"48",x"d0",x"ff",x"78"),
   228 => (x"ff",x"78",x"c3",x"c4"),
   229 => (x"ff",x"c3",x"48",x"d4"),
   230 => (x"c0",x"1e",x"72",x"78"),
   231 => (x"d1",x"c1",x"f0",x"ff"),
   232 => (x"87",x"ef",x"f5",x"49"),
   233 => (x"98",x"70",x"86",x"c4"),
   234 => (x"c8",x"87",x"d2",x"05"),
   235 => (x"66",x"cc",x"1e",x"c0"),
   236 => (x"87",x"e6",x"fd",x"49"),
   237 => (x"4b",x"70",x"86",x"c4"),
   238 => (x"c2",x"48",x"d0",x"ff"),
   239 => (x"f5",x"48",x"73",x"78"),
   240 => (x"5e",x"0e",x"87",x"cd"),
   241 => (x"0e",x"5d",x"5c",x"5b"),
   242 => (x"ff",x"c0",x"1e",x"c0"),
   243 => (x"49",x"c9",x"c1",x"f0"),
   244 => (x"d2",x"87",x"c0",x"f5"),
   245 => (x"f8",x"ce",x"c2",x"1e"),
   246 => (x"87",x"fe",x"fc",x"49"),
   247 => (x"4c",x"c0",x"86",x"c8"),
   248 => (x"b7",x"d2",x"84",x"c1"),
   249 => (x"87",x"f8",x"04",x"ac"),
   250 => (x"97",x"f8",x"ce",x"c2"),
   251 => (x"c0",x"c3",x"49",x"bf"),
   252 => (x"a9",x"c0",x"c1",x"99"),
   253 => (x"87",x"e7",x"c0",x"05"),
   254 => (x"97",x"ff",x"ce",x"c2"),
   255 => (x"31",x"d0",x"49",x"bf"),
   256 => (x"97",x"c0",x"cf",x"c2"),
   257 => (x"32",x"c8",x"4a",x"bf"),
   258 => (x"cf",x"c2",x"b1",x"72"),
   259 => (x"4a",x"bf",x"97",x"c1"),
   260 => (x"cf",x"4c",x"71",x"b1"),
   261 => (x"9c",x"ff",x"ff",x"ff"),
   262 => (x"34",x"ca",x"84",x"c1"),
   263 => (x"c2",x"87",x"e7",x"c1"),
   264 => (x"bf",x"97",x"c1",x"cf"),
   265 => (x"c6",x"31",x"c1",x"49"),
   266 => (x"c2",x"cf",x"c2",x"99"),
   267 => (x"c7",x"4a",x"bf",x"97"),
   268 => (x"b1",x"72",x"2a",x"b7"),
   269 => (x"97",x"fd",x"ce",x"c2"),
   270 => (x"cf",x"4d",x"4a",x"bf"),
   271 => (x"fe",x"ce",x"c2",x"9d"),
   272 => (x"c3",x"4a",x"bf",x"97"),
   273 => (x"c2",x"32",x"ca",x"9a"),
   274 => (x"bf",x"97",x"ff",x"ce"),
   275 => (x"73",x"33",x"c2",x"4b"),
   276 => (x"c0",x"cf",x"c2",x"b2"),
   277 => (x"c3",x"4b",x"bf",x"97"),
   278 => (x"b7",x"c6",x"9b",x"c0"),
   279 => (x"c2",x"b2",x"73",x"2b"),
   280 => (x"71",x"48",x"c1",x"81"),
   281 => (x"c1",x"49",x"70",x"30"),
   282 => (x"70",x"30",x"75",x"48"),
   283 => (x"c1",x"4c",x"72",x"4d"),
   284 => (x"c8",x"94",x"71",x"84"),
   285 => (x"06",x"ad",x"b7",x"c0"),
   286 => (x"34",x"c1",x"87",x"cc"),
   287 => (x"c0",x"c8",x"2d",x"b7"),
   288 => (x"ff",x"01",x"ad",x"b7"),
   289 => (x"48",x"74",x"87",x"f4"),
   290 => (x"0e",x"87",x"c0",x"f2"),
   291 => (x"5d",x"5c",x"5b",x"5e"),
   292 => (x"c2",x"86",x"f8",x"0e"),
   293 => (x"c0",x"48",x"de",x"d7"),
   294 => (x"d6",x"cf",x"c2",x"78"),
   295 => (x"fb",x"49",x"c0",x"1e"),
   296 => (x"86",x"c4",x"87",x"de"),
   297 => (x"c5",x"05",x"98",x"70"),
   298 => (x"c9",x"48",x"c0",x"87"),
   299 => (x"4d",x"c0",x"87",x"ce"),
   300 => (x"ed",x"c0",x"7e",x"c1"),
   301 => (x"c2",x"49",x"bf",x"f3"),
   302 => (x"71",x"4a",x"cc",x"d0"),
   303 => (x"e9",x"ee",x"4b",x"c8"),
   304 => (x"05",x"98",x"70",x"87"),
   305 => (x"7e",x"c0",x"87",x"c2"),
   306 => (x"bf",x"ef",x"ed",x"c0"),
   307 => (x"e8",x"d0",x"c2",x"49"),
   308 => (x"4b",x"c8",x"71",x"4a"),
   309 => (x"70",x"87",x"d3",x"ee"),
   310 => (x"87",x"c2",x"05",x"98"),
   311 => (x"02",x"6e",x"7e",x"c0"),
   312 => (x"c2",x"87",x"fd",x"c0"),
   313 => (x"4d",x"bf",x"dc",x"d6"),
   314 => (x"9f",x"d4",x"d7",x"c2"),
   315 => (x"c5",x"48",x"7e",x"bf"),
   316 => (x"05",x"a8",x"ea",x"d6"),
   317 => (x"d6",x"c2",x"87",x"c7"),
   318 => (x"ce",x"4d",x"bf",x"dc"),
   319 => (x"ca",x"48",x"6e",x"87"),
   320 => (x"02",x"a8",x"d5",x"e9"),
   321 => (x"48",x"c0",x"87",x"c5"),
   322 => (x"c2",x"87",x"f1",x"c7"),
   323 => (x"75",x"1e",x"d6",x"cf"),
   324 => (x"87",x"ec",x"f9",x"49"),
   325 => (x"98",x"70",x"86",x"c4"),
   326 => (x"c0",x"87",x"c5",x"05"),
   327 => (x"87",x"dc",x"c7",x"48"),
   328 => (x"bf",x"ef",x"ed",x"c0"),
   329 => (x"e8",x"d0",x"c2",x"49"),
   330 => (x"4b",x"c8",x"71",x"4a"),
   331 => (x"70",x"87",x"fb",x"ec"),
   332 => (x"87",x"c8",x"05",x"98"),
   333 => (x"48",x"de",x"d7",x"c2"),
   334 => (x"87",x"da",x"78",x"c1"),
   335 => (x"bf",x"f3",x"ed",x"c0"),
   336 => (x"cc",x"d0",x"c2",x"49"),
   337 => (x"4b",x"c8",x"71",x"4a"),
   338 => (x"70",x"87",x"df",x"ec"),
   339 => (x"c5",x"c0",x"02",x"98"),
   340 => (x"c6",x"48",x"c0",x"87"),
   341 => (x"d7",x"c2",x"87",x"e6"),
   342 => (x"49",x"bf",x"97",x"d4"),
   343 => (x"05",x"a9",x"d5",x"c1"),
   344 => (x"c2",x"87",x"cd",x"c0"),
   345 => (x"bf",x"97",x"d5",x"d7"),
   346 => (x"a9",x"ea",x"c2",x"49"),
   347 => (x"87",x"c5",x"c0",x"02"),
   348 => (x"c7",x"c6",x"48",x"c0"),
   349 => (x"d6",x"cf",x"c2",x"87"),
   350 => (x"48",x"7e",x"bf",x"97"),
   351 => (x"02",x"a8",x"e9",x"c3"),
   352 => (x"6e",x"87",x"ce",x"c0"),
   353 => (x"a8",x"eb",x"c3",x"48"),
   354 => (x"87",x"c5",x"c0",x"02"),
   355 => (x"eb",x"c5",x"48",x"c0"),
   356 => (x"e1",x"cf",x"c2",x"87"),
   357 => (x"99",x"49",x"bf",x"97"),
   358 => (x"87",x"cc",x"c0",x"05"),
   359 => (x"97",x"e2",x"cf",x"c2"),
   360 => (x"a9",x"c2",x"49",x"bf"),
   361 => (x"87",x"c5",x"c0",x"02"),
   362 => (x"cf",x"c5",x"48",x"c0"),
   363 => (x"e3",x"cf",x"c2",x"87"),
   364 => (x"c2",x"48",x"bf",x"97"),
   365 => (x"70",x"58",x"da",x"d7"),
   366 => (x"88",x"c1",x"48",x"4c"),
   367 => (x"58",x"de",x"d7",x"c2"),
   368 => (x"97",x"e4",x"cf",x"c2"),
   369 => (x"81",x"75",x"49",x"bf"),
   370 => (x"97",x"e5",x"cf",x"c2"),
   371 => (x"32",x"c8",x"4a",x"bf"),
   372 => (x"c2",x"7e",x"a1",x"72"),
   373 => (x"6e",x"48",x"eb",x"db"),
   374 => (x"e6",x"cf",x"c2",x"78"),
   375 => (x"c8",x"48",x"bf",x"97"),
   376 => (x"d7",x"c2",x"58",x"a6"),
   377 => (x"c2",x"02",x"bf",x"de"),
   378 => (x"ed",x"c0",x"87",x"d4"),
   379 => (x"c2",x"49",x"bf",x"ef"),
   380 => (x"71",x"4a",x"e8",x"d0"),
   381 => (x"f1",x"e9",x"4b",x"c8"),
   382 => (x"02",x"98",x"70",x"87"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f8",x"c3",x"48"),
   385 => (x"bf",x"d6",x"d7",x"c2"),
   386 => (x"ff",x"db",x"c2",x"4c"),
   387 => (x"fb",x"cf",x"c2",x"5c"),
   388 => (x"c8",x"49",x"bf",x"97"),
   389 => (x"fa",x"cf",x"c2",x"31"),
   390 => (x"a1",x"4a",x"bf",x"97"),
   391 => (x"fc",x"cf",x"c2",x"49"),
   392 => (x"d0",x"4a",x"bf",x"97"),
   393 => (x"49",x"a1",x"72",x"32"),
   394 => (x"97",x"fd",x"cf",x"c2"),
   395 => (x"32",x"d8",x"4a",x"bf"),
   396 => (x"c4",x"49",x"a1",x"72"),
   397 => (x"db",x"c2",x"91",x"66"),
   398 => (x"c2",x"81",x"bf",x"eb"),
   399 => (x"c2",x"59",x"f3",x"db"),
   400 => (x"bf",x"97",x"c3",x"d0"),
   401 => (x"c2",x"32",x"c8",x"4a"),
   402 => (x"bf",x"97",x"c2",x"d0"),
   403 => (x"c2",x"4a",x"a2",x"4b"),
   404 => (x"bf",x"97",x"c4",x"d0"),
   405 => (x"73",x"33",x"d0",x"4b"),
   406 => (x"d0",x"c2",x"4a",x"a2"),
   407 => (x"4b",x"bf",x"97",x"c5"),
   408 => (x"33",x"d8",x"9b",x"cf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"c2",x"5a",x"f7",x"db"),
   411 => (x"4a",x"bf",x"f3",x"db"),
   412 => (x"92",x"74",x"8a",x"c2"),
   413 => (x"48",x"f7",x"db",x"c2"),
   414 => (x"c1",x"78",x"a1",x"72"),
   415 => (x"cf",x"c2",x"87",x"ca"),
   416 => (x"49",x"bf",x"97",x"e8"),
   417 => (x"cf",x"c2",x"31",x"c8"),
   418 => (x"4a",x"bf",x"97",x"e7"),
   419 => (x"d7",x"c2",x"49",x"a1"),
   420 => (x"d7",x"c2",x"59",x"e6"),
   421 => (x"c5",x"49",x"bf",x"e2"),
   422 => (x"81",x"ff",x"c7",x"31"),
   423 => (x"db",x"c2",x"29",x"c9"),
   424 => (x"cf",x"c2",x"59",x"ff"),
   425 => (x"4a",x"bf",x"97",x"ed"),
   426 => (x"cf",x"c2",x"32",x"c8"),
   427 => (x"4b",x"bf",x"97",x"ec"),
   428 => (x"66",x"c4",x"4a",x"a2"),
   429 => (x"c2",x"82",x"6e",x"92"),
   430 => (x"c2",x"5a",x"fb",x"db"),
   431 => (x"c0",x"48",x"f3",x"db"),
   432 => (x"ef",x"db",x"c2",x"78"),
   433 => (x"78",x"a1",x"72",x"48"),
   434 => (x"48",x"ff",x"db",x"c2"),
   435 => (x"bf",x"f3",x"db",x"c2"),
   436 => (x"c3",x"dc",x"c2",x"78"),
   437 => (x"f7",x"db",x"c2",x"48"),
   438 => (x"d7",x"c2",x"78",x"bf"),
   439 => (x"c0",x"02",x"bf",x"de"),
   440 => (x"48",x"74",x"87",x"c9"),
   441 => (x"7e",x"70",x"30",x"c4"),
   442 => (x"c2",x"87",x"c9",x"c0"),
   443 => (x"48",x"bf",x"fb",x"db"),
   444 => (x"7e",x"70",x"30",x"c4"),
   445 => (x"48",x"e2",x"d7",x"c2"),
   446 => (x"48",x"c1",x"78",x"6e"),
   447 => (x"4d",x"26",x"8e",x"f8"),
   448 => (x"4b",x"26",x"4c",x"26"),
   449 => (x"5e",x"0e",x"4f",x"26"),
   450 => (x"0e",x"5d",x"5c",x"5b"),
   451 => (x"d7",x"c2",x"4a",x"71"),
   452 => (x"cb",x"02",x"bf",x"de"),
   453 => (x"c7",x"4b",x"72",x"87"),
   454 => (x"c1",x"4c",x"72",x"2b"),
   455 => (x"87",x"c9",x"9c",x"ff"),
   456 => (x"2b",x"c8",x"4b",x"72"),
   457 => (x"ff",x"c3",x"4c",x"72"),
   458 => (x"eb",x"db",x"c2",x"9c"),
   459 => (x"ed",x"c0",x"83",x"bf"),
   460 => (x"02",x"ab",x"bf",x"eb"),
   461 => (x"ed",x"c0",x"87",x"d9"),
   462 => (x"cf",x"c2",x"5b",x"ef"),
   463 => (x"49",x"73",x"1e",x"d6"),
   464 => (x"c4",x"87",x"fd",x"f0"),
   465 => (x"05",x"98",x"70",x"86"),
   466 => (x"48",x"c0",x"87",x"c5"),
   467 => (x"c2",x"87",x"e6",x"c0"),
   468 => (x"02",x"bf",x"de",x"d7"),
   469 => (x"49",x"74",x"87",x"d2"),
   470 => (x"cf",x"c2",x"91",x"c4"),
   471 => (x"4d",x"69",x"81",x"d6"),
   472 => (x"ff",x"ff",x"ff",x"cf"),
   473 => (x"87",x"cb",x"9d",x"ff"),
   474 => (x"91",x"c2",x"49",x"74"),
   475 => (x"81",x"d6",x"cf",x"c2"),
   476 => (x"75",x"4d",x"69",x"9f"),
   477 => (x"87",x"c6",x"fe",x"48"),
   478 => (x"5c",x"5b",x"5e",x"0e"),
   479 => (x"86",x"f8",x"0e",x"5d"),
   480 => (x"05",x"9c",x"4c",x"71"),
   481 => (x"48",x"c0",x"87",x"c5"),
   482 => (x"c8",x"87",x"c1",x"c3"),
   483 => (x"48",x"6e",x"7e",x"a4"),
   484 => (x"66",x"d8",x"78",x"c0"),
   485 => (x"d8",x"87",x"c7",x"02"),
   486 => (x"05",x"bf",x"97",x"66"),
   487 => (x"48",x"c0",x"87",x"c5"),
   488 => (x"c0",x"87",x"e9",x"c2"),
   489 => (x"c7",x"49",x"c1",x"1e"),
   490 => (x"86",x"c4",x"87",x"e6"),
   491 => (x"02",x"9d",x"4d",x"70"),
   492 => (x"c2",x"87",x"c2",x"c1"),
   493 => (x"d8",x"4a",x"e6",x"d7"),
   494 => (x"d2",x"e2",x"49",x"66"),
   495 => (x"02",x"98",x"70",x"87"),
   496 => (x"75",x"87",x"f2",x"c0"),
   497 => (x"49",x"66",x"d8",x"4a"),
   498 => (x"f7",x"e2",x"4b",x"cb"),
   499 => (x"02",x"98",x"70",x"87"),
   500 => (x"c0",x"87",x"e2",x"c0"),
   501 => (x"02",x"9d",x"75",x"1e"),
   502 => (x"a6",x"c8",x"87",x"c7"),
   503 => (x"c5",x"78",x"c0",x"48"),
   504 => (x"48",x"a6",x"c8",x"87"),
   505 => (x"66",x"c8",x"78",x"c1"),
   506 => (x"87",x"e4",x"c6",x"49"),
   507 => (x"4d",x"70",x"86",x"c4"),
   508 => (x"fe",x"fe",x"05",x"9d"),
   509 => (x"02",x"9d",x"75",x"87"),
   510 => (x"dc",x"87",x"cf",x"c1"),
   511 => (x"48",x"6e",x"49",x"a5"),
   512 => (x"a5",x"da",x"78",x"69"),
   513 => (x"48",x"a6",x"c4",x"49"),
   514 => (x"9f",x"78",x"a4",x"c4"),
   515 => (x"66",x"c4",x"48",x"69"),
   516 => (x"d7",x"c2",x"78",x"08"),
   517 => (x"d2",x"02",x"bf",x"de"),
   518 => (x"49",x"a5",x"d4",x"87"),
   519 => (x"c0",x"49",x"69",x"9f"),
   520 => (x"71",x"99",x"ff",x"ff"),
   521 => (x"70",x"30",x"d0",x"48"),
   522 => (x"c0",x"87",x"c2",x"7e"),
   523 => (x"48",x"49",x"6e",x"7e"),
   524 => (x"80",x"bf",x"66",x"c4"),
   525 => (x"78",x"08",x"66",x"c4"),
   526 => (x"a4",x"cc",x"7c",x"c0"),
   527 => (x"bf",x"66",x"c4",x"49"),
   528 => (x"49",x"a4",x"d0",x"79"),
   529 => (x"48",x"c1",x"79",x"c0"),
   530 => (x"48",x"c0",x"87",x"c2"),
   531 => (x"ed",x"fa",x"8e",x"f8"),
   532 => (x"5b",x"5e",x"0e",x"87"),
   533 => (x"71",x"0e",x"5d",x"5c"),
   534 => (x"c1",x"02",x"9c",x"4c"),
   535 => (x"a4",x"c8",x"87",x"ca"),
   536 => (x"c1",x"02",x"69",x"49"),
   537 => (x"66",x"d0",x"87",x"c2"),
   538 => (x"82",x"49",x"6c",x"4a"),
   539 => (x"d0",x"5a",x"a6",x"d4"),
   540 => (x"c2",x"b9",x"4d",x"66"),
   541 => (x"4a",x"bf",x"da",x"d7"),
   542 => (x"99",x"72",x"ba",x"ff"),
   543 => (x"c0",x"02",x"99",x"71"),
   544 => (x"a4",x"c4",x"87",x"e4"),
   545 => (x"f9",x"49",x"6b",x"4b"),
   546 => (x"7b",x"70",x"87",x"fc"),
   547 => (x"bf",x"d6",x"d7",x"c2"),
   548 => (x"71",x"81",x"6c",x"49"),
   549 => (x"c2",x"b9",x"75",x"7c"),
   550 => (x"4a",x"bf",x"da",x"d7"),
   551 => (x"99",x"72",x"ba",x"ff"),
   552 => (x"ff",x"05",x"99",x"71"),
   553 => (x"7c",x"75",x"87",x"dc"),
   554 => (x"1e",x"87",x"d3",x"f9"),
   555 => (x"4b",x"71",x"1e",x"73"),
   556 => (x"87",x"c7",x"02",x"9b"),
   557 => (x"69",x"49",x"a3",x"c8"),
   558 => (x"c0",x"87",x"c5",x"05"),
   559 => (x"87",x"f7",x"c0",x"48"),
   560 => (x"bf",x"ef",x"db",x"c2"),
   561 => (x"49",x"a3",x"c4",x"4a"),
   562 => (x"89",x"c2",x"49",x"69"),
   563 => (x"bf",x"d6",x"d7",x"c2"),
   564 => (x"4a",x"a2",x"71",x"91"),
   565 => (x"bf",x"da",x"d7",x"c2"),
   566 => (x"71",x"99",x"6b",x"49"),
   567 => (x"ed",x"c0",x"4a",x"a2"),
   568 => (x"66",x"c8",x"5a",x"ef"),
   569 => (x"ea",x"49",x"72",x"1e"),
   570 => (x"86",x"c4",x"87",x"d6"),
   571 => (x"c4",x"05",x"98",x"70"),
   572 => (x"c2",x"48",x"c0",x"87"),
   573 => (x"f8",x"48",x"c1",x"87"),
   574 => (x"73",x"1e",x"87",x"c8"),
   575 => (x"9b",x"4b",x"71",x"1e"),
   576 => (x"87",x"e4",x"c0",x"02"),
   577 => (x"5b",x"c3",x"dc",x"c2"),
   578 => (x"8a",x"c2",x"4a",x"73"),
   579 => (x"bf",x"d6",x"d7",x"c2"),
   580 => (x"db",x"c2",x"92",x"49"),
   581 => (x"72",x"48",x"bf",x"ef"),
   582 => (x"c7",x"dc",x"c2",x"80"),
   583 => (x"c4",x"48",x"71",x"58"),
   584 => (x"e6",x"d7",x"c2",x"30"),
   585 => (x"87",x"ed",x"c0",x"58"),
   586 => (x"48",x"ff",x"db",x"c2"),
   587 => (x"bf",x"f3",x"db",x"c2"),
   588 => (x"c3",x"dc",x"c2",x"78"),
   589 => (x"f7",x"db",x"c2",x"48"),
   590 => (x"d7",x"c2",x"78",x"bf"),
   591 => (x"c9",x"02",x"bf",x"de"),
   592 => (x"d6",x"d7",x"c2",x"87"),
   593 => (x"31",x"c4",x"49",x"bf"),
   594 => (x"db",x"c2",x"87",x"c7"),
   595 => (x"c4",x"49",x"bf",x"fb"),
   596 => (x"e6",x"d7",x"c2",x"31"),
   597 => (x"87",x"ea",x"f6",x"59"),
   598 => (x"5c",x"5b",x"5e",x"0e"),
   599 => (x"c0",x"4a",x"71",x"0e"),
   600 => (x"02",x"9a",x"72",x"4b"),
   601 => (x"da",x"87",x"e1",x"c0"),
   602 => (x"69",x"9f",x"49",x"a2"),
   603 => (x"de",x"d7",x"c2",x"4b"),
   604 => (x"87",x"cf",x"02",x"bf"),
   605 => (x"9f",x"49",x"a2",x"d4"),
   606 => (x"c0",x"4c",x"49",x"69"),
   607 => (x"d0",x"9c",x"ff",x"ff"),
   608 => (x"c0",x"87",x"c2",x"34"),
   609 => (x"b3",x"49",x"74",x"4c"),
   610 => (x"ed",x"fd",x"49",x"73"),
   611 => (x"87",x"f0",x"f5",x"87"),
   612 => (x"5c",x"5b",x"5e",x"0e"),
   613 => (x"86",x"f4",x"0e",x"5d"),
   614 => (x"7e",x"c0",x"4a",x"71"),
   615 => (x"d8",x"02",x"9a",x"72"),
   616 => (x"d2",x"cf",x"c2",x"87"),
   617 => (x"c2",x"78",x"c0",x"48"),
   618 => (x"c2",x"48",x"ca",x"cf"),
   619 => (x"78",x"bf",x"c3",x"dc"),
   620 => (x"48",x"ce",x"cf",x"c2"),
   621 => (x"bf",x"ff",x"db",x"c2"),
   622 => (x"f3",x"d7",x"c2",x"78"),
   623 => (x"c2",x"50",x"c0",x"48"),
   624 => (x"49",x"bf",x"e2",x"d7"),
   625 => (x"bf",x"d2",x"cf",x"c2"),
   626 => (x"03",x"aa",x"71",x"4a"),
   627 => (x"72",x"87",x"c9",x"c4"),
   628 => (x"05",x"99",x"cf",x"49"),
   629 => (x"c0",x"87",x"e9",x"c0"),
   630 => (x"c2",x"48",x"eb",x"ed"),
   631 => (x"78",x"bf",x"ca",x"cf"),
   632 => (x"1e",x"d6",x"cf",x"c2"),
   633 => (x"bf",x"ca",x"cf",x"c2"),
   634 => (x"ca",x"cf",x"c2",x"49"),
   635 => (x"78",x"a1",x"c1",x"48"),
   636 => (x"87",x"cc",x"e6",x"71"),
   637 => (x"ed",x"c0",x"86",x"c4"),
   638 => (x"cf",x"c2",x"48",x"e7"),
   639 => (x"87",x"cc",x"78",x"d6"),
   640 => (x"bf",x"e7",x"ed",x"c0"),
   641 => (x"80",x"e0",x"c0",x"48"),
   642 => (x"58",x"eb",x"ed",x"c0"),
   643 => (x"bf",x"d2",x"cf",x"c2"),
   644 => (x"c2",x"80",x"c1",x"48"),
   645 => (x"27",x"58",x"d6",x"cf"),
   646 => (x"00",x"00",x"0b",x"67"),
   647 => (x"4d",x"bf",x"97",x"bf"),
   648 => (x"e3",x"c2",x"02",x"9d"),
   649 => (x"ad",x"e5",x"c3",x"87"),
   650 => (x"87",x"dc",x"c2",x"02"),
   651 => (x"bf",x"e7",x"ed",x"c0"),
   652 => (x"49",x"a3",x"cb",x"4b"),
   653 => (x"ac",x"cf",x"4c",x"11"),
   654 => (x"87",x"d2",x"c1",x"05"),
   655 => (x"99",x"df",x"49",x"75"),
   656 => (x"91",x"cd",x"89",x"c1"),
   657 => (x"81",x"e6",x"d7",x"c2"),
   658 => (x"12",x"4a",x"a3",x"c1"),
   659 => (x"4a",x"a3",x"c3",x"51"),
   660 => (x"a3",x"c5",x"51",x"12"),
   661 => (x"c7",x"51",x"12",x"4a"),
   662 => (x"51",x"12",x"4a",x"a3"),
   663 => (x"12",x"4a",x"a3",x"c9"),
   664 => (x"4a",x"a3",x"ce",x"51"),
   665 => (x"a3",x"d0",x"51",x"12"),
   666 => (x"d2",x"51",x"12",x"4a"),
   667 => (x"51",x"12",x"4a",x"a3"),
   668 => (x"12",x"4a",x"a3",x"d4"),
   669 => (x"4a",x"a3",x"d6",x"51"),
   670 => (x"a3",x"d8",x"51",x"12"),
   671 => (x"dc",x"51",x"12",x"4a"),
   672 => (x"51",x"12",x"4a",x"a3"),
   673 => (x"12",x"4a",x"a3",x"de"),
   674 => (x"c0",x"7e",x"c1",x"51"),
   675 => (x"49",x"74",x"87",x"fa"),
   676 => (x"c0",x"05",x"99",x"c8"),
   677 => (x"49",x"74",x"87",x"eb"),
   678 => (x"d1",x"05",x"99",x"d0"),
   679 => (x"02",x"66",x"dc",x"87"),
   680 => (x"73",x"87",x"cb",x"c0"),
   681 => (x"0f",x"66",x"dc",x"49"),
   682 => (x"c0",x"02",x"98",x"70"),
   683 => (x"05",x"6e",x"87",x"d3"),
   684 => (x"c2",x"87",x"c6",x"c0"),
   685 => (x"c0",x"48",x"e6",x"d7"),
   686 => (x"e7",x"ed",x"c0",x"50"),
   687 => (x"e1",x"c2",x"48",x"bf"),
   688 => (x"f3",x"d7",x"c2",x"87"),
   689 => (x"7e",x"50",x"c0",x"48"),
   690 => (x"bf",x"e2",x"d7",x"c2"),
   691 => (x"d2",x"cf",x"c2",x"49"),
   692 => (x"aa",x"71",x"4a",x"bf"),
   693 => (x"87",x"f7",x"fb",x"04"),
   694 => (x"bf",x"c3",x"dc",x"c2"),
   695 => (x"87",x"c8",x"c0",x"05"),
   696 => (x"bf",x"de",x"d7",x"c2"),
   697 => (x"87",x"f8",x"c1",x"02"),
   698 => (x"bf",x"ce",x"cf",x"c2"),
   699 => (x"87",x"d6",x"f0",x"49"),
   700 => (x"cf",x"c2",x"49",x"70"),
   701 => (x"a6",x"c4",x"59",x"d2"),
   702 => (x"ce",x"cf",x"c2",x"48"),
   703 => (x"d7",x"c2",x"78",x"bf"),
   704 => (x"c0",x"02",x"bf",x"de"),
   705 => (x"66",x"c4",x"87",x"d8"),
   706 => (x"ff",x"ff",x"cf",x"49"),
   707 => (x"a9",x"99",x"f8",x"ff"),
   708 => (x"87",x"c5",x"c0",x"02"),
   709 => (x"e1",x"c0",x"4c",x"c0"),
   710 => (x"c0",x"4c",x"c1",x"87"),
   711 => (x"66",x"c4",x"87",x"dc"),
   712 => (x"f8",x"ff",x"cf",x"49"),
   713 => (x"c0",x"02",x"a9",x"99"),
   714 => (x"a6",x"c8",x"87",x"c8"),
   715 => (x"c0",x"78",x"c0",x"48"),
   716 => (x"a6",x"c8",x"87",x"c5"),
   717 => (x"c8",x"78",x"c1",x"48"),
   718 => (x"9c",x"74",x"4c",x"66"),
   719 => (x"87",x"e0",x"c0",x"05"),
   720 => (x"c2",x"49",x"66",x"c4"),
   721 => (x"d6",x"d7",x"c2",x"89"),
   722 => (x"c2",x"91",x"4a",x"bf"),
   723 => (x"4a",x"bf",x"ef",x"db"),
   724 => (x"48",x"ca",x"cf",x"c2"),
   725 => (x"c2",x"78",x"a1",x"72"),
   726 => (x"c0",x"48",x"d2",x"cf"),
   727 => (x"87",x"df",x"f9",x"78"),
   728 => (x"8e",x"f4",x"48",x"c0"),
   729 => (x"00",x"87",x"d7",x"ee"),
   730 => (x"ff",x"00",x"00",x"00"),
   731 => (x"77",x"ff",x"ff",x"ff"),
   732 => (x"80",x"00",x"00",x"0b"),
   733 => (x"46",x"00",x"00",x"0b"),
   734 => (x"32",x"33",x"54",x"41"),
   735 => (x"00",x"20",x"20",x"20"),
   736 => (x"31",x"54",x"41",x"46"),
   737 => (x"20",x"20",x"20",x"36"),
   738 => (x"d4",x"ff",x"1e",x"00"),
   739 => (x"78",x"ff",x"c3",x"48"),
   740 => (x"4f",x"26",x"48",x"68"),
   741 => (x"48",x"d4",x"ff",x"1e"),
   742 => (x"ff",x"78",x"ff",x"c3"),
   743 => (x"e1",x"c0",x"48",x"d0"),
   744 => (x"48",x"d4",x"ff",x"78"),
   745 => (x"dc",x"c2",x"78",x"d4"),
   746 => (x"d4",x"ff",x"48",x"c7"),
   747 => (x"4f",x"26",x"50",x"bf"),
   748 => (x"48",x"d0",x"ff",x"1e"),
   749 => (x"26",x"78",x"e0",x"c0"),
   750 => (x"cc",x"ff",x"1e",x"4f"),
   751 => (x"99",x"49",x"70",x"87"),
   752 => (x"c0",x"87",x"c6",x"02"),
   753 => (x"f1",x"05",x"a9",x"fb"),
   754 => (x"26",x"48",x"71",x"87"),
   755 => (x"5b",x"5e",x"0e",x"4f"),
   756 => (x"4b",x"71",x"0e",x"5c"),
   757 => (x"f0",x"fe",x"4c",x"c0"),
   758 => (x"99",x"49",x"70",x"87"),
   759 => (x"87",x"f9",x"c0",x"02"),
   760 => (x"02",x"a9",x"ec",x"c0"),
   761 => (x"c0",x"87",x"f2",x"c0"),
   762 => (x"c0",x"02",x"a9",x"fb"),
   763 => (x"66",x"cc",x"87",x"eb"),
   764 => (x"c7",x"03",x"ac",x"b7"),
   765 => (x"02",x"66",x"d0",x"87"),
   766 => (x"53",x"71",x"87",x"c2"),
   767 => (x"c2",x"02",x"99",x"71"),
   768 => (x"fe",x"84",x"c1",x"87"),
   769 => (x"49",x"70",x"87",x"c3"),
   770 => (x"87",x"cd",x"02",x"99"),
   771 => (x"02",x"a9",x"ec",x"c0"),
   772 => (x"fb",x"c0",x"87",x"c7"),
   773 => (x"d5",x"ff",x"05",x"a9"),
   774 => (x"02",x"66",x"d0",x"87"),
   775 => (x"97",x"c0",x"87",x"c3"),
   776 => (x"a9",x"ec",x"c0",x"7b"),
   777 => (x"74",x"87",x"c4",x"05"),
   778 => (x"74",x"87",x"c5",x"4a"),
   779 => (x"8a",x"0a",x"c0",x"4a"),
   780 => (x"87",x"c2",x"48",x"72"),
   781 => (x"4c",x"26",x"4d",x"26"),
   782 => (x"4f",x"26",x"4b",x"26"),
   783 => (x"87",x"c9",x"fd",x"1e"),
   784 => (x"c0",x"4a",x"49",x"70"),
   785 => (x"c9",x"04",x"aa",x"f0"),
   786 => (x"aa",x"f9",x"c0",x"87"),
   787 => (x"c0",x"87",x"c3",x"01"),
   788 => (x"c1",x"c1",x"8a",x"f0"),
   789 => (x"87",x"c9",x"04",x"aa"),
   790 => (x"01",x"aa",x"da",x"c1"),
   791 => (x"f7",x"c0",x"87",x"c3"),
   792 => (x"26",x"48",x"72",x"8a"),
   793 => (x"5b",x"5e",x"0e",x"4f"),
   794 => (x"f8",x"0e",x"5d",x"5c"),
   795 => (x"c0",x"4c",x"71",x"86"),
   796 => (x"87",x"e0",x"fc",x"4d"),
   797 => (x"f4",x"c0",x"4b",x"c0"),
   798 => (x"49",x"bf",x"97",x"c4"),
   799 => (x"cf",x"04",x"a9",x"c0"),
   800 => (x"87",x"f5",x"fc",x"87"),
   801 => (x"f4",x"c0",x"83",x"c1"),
   802 => (x"49",x"bf",x"97",x"c4"),
   803 => (x"87",x"f1",x"06",x"ab"),
   804 => (x"97",x"c4",x"f4",x"c0"),
   805 => (x"87",x"cf",x"02",x"bf"),
   806 => (x"70",x"87",x"ee",x"fb"),
   807 => (x"c6",x"02",x"99",x"49"),
   808 => (x"a9",x"ec",x"c0",x"87"),
   809 => (x"c0",x"87",x"f1",x"05"),
   810 => (x"87",x"dd",x"fb",x"4b"),
   811 => (x"d8",x"fb",x"7e",x"70"),
   812 => (x"58",x"a6",x"c8",x"87"),
   813 => (x"70",x"87",x"d2",x"fb"),
   814 => (x"c8",x"83",x"c1",x"4a"),
   815 => (x"69",x"97",x"49",x"a4"),
   816 => (x"05",x"a9",x"6e",x"49"),
   817 => (x"a4",x"c9",x"87",x"da"),
   818 => (x"49",x"69",x"97",x"49"),
   819 => (x"05",x"a9",x"66",x"c4"),
   820 => (x"a4",x"ca",x"87",x"ce"),
   821 => (x"49",x"69",x"97",x"49"),
   822 => (x"87",x"c4",x"05",x"aa"),
   823 => (x"87",x"d4",x"4d",x"c1"),
   824 => (x"ec",x"c0",x"48",x"6e"),
   825 => (x"87",x"c8",x"02",x"a8"),
   826 => (x"fb",x"c0",x"48",x"6e"),
   827 => (x"87",x"c4",x"05",x"a8"),
   828 => (x"4d",x"c1",x"4b",x"c0"),
   829 => (x"fe",x"02",x"9d",x"75"),
   830 => (x"f3",x"fa",x"87",x"ef"),
   831 => (x"f8",x"48",x"73",x"87"),
   832 => (x"87",x"f0",x"fc",x"8e"),
   833 => (x"5b",x"5e",x"0e",x"00"),
   834 => (x"f8",x"0e",x"5d",x"5c"),
   835 => (x"ff",x"7e",x"71",x"86"),
   836 => (x"1e",x"6e",x"4b",x"d4"),
   837 => (x"49",x"cc",x"dc",x"c2"),
   838 => (x"c4",x"87",x"dd",x"e9"),
   839 => (x"02",x"98",x"70",x"86"),
   840 => (x"c1",x"87",x"ec",x"c4"),
   841 => (x"4d",x"bf",x"df",x"de"),
   842 => (x"f8",x"fc",x"49",x"6e"),
   843 => (x"58",x"a6",x"c8",x"87"),
   844 => (x"c5",x"05",x"98",x"70"),
   845 => (x"48",x"a6",x"c4",x"87"),
   846 => (x"d0",x"ff",x"78",x"c1"),
   847 => (x"c1",x"78",x"c5",x"48"),
   848 => (x"66",x"c4",x"7b",x"d5"),
   849 => (x"c6",x"89",x"c1",x"49"),
   850 => (x"dd",x"de",x"c1",x"31"),
   851 => (x"48",x"4a",x"bf",x"97"),
   852 => (x"7b",x"70",x"b0",x"71"),
   853 => (x"c4",x"48",x"d0",x"ff"),
   854 => (x"c7",x"dc",x"c2",x"78"),
   855 => (x"d0",x"49",x"bf",x"97"),
   856 => (x"87",x"d7",x"02",x"99"),
   857 => (x"d6",x"c1",x"78",x"c5"),
   858 => (x"c3",x"4a",x"c0",x"7b"),
   859 => (x"82",x"c1",x"7b",x"ff"),
   860 => (x"04",x"aa",x"e0",x"c0"),
   861 => (x"d0",x"ff",x"87",x"f5"),
   862 => (x"c3",x"78",x"c4",x"48"),
   863 => (x"d0",x"ff",x"7b",x"ff"),
   864 => (x"c1",x"78",x"c5",x"48"),
   865 => (x"7b",x"c1",x"7b",x"d3"),
   866 => (x"b7",x"c0",x"78",x"c4"),
   867 => (x"ed",x"c2",x"06",x"ad"),
   868 => (x"d4",x"dc",x"c2",x"87"),
   869 => (x"9c",x"8d",x"4c",x"bf"),
   870 => (x"87",x"c4",x"c2",x"02"),
   871 => (x"7e",x"d6",x"cf",x"c2"),
   872 => (x"c8",x"48",x"a6",x"c4"),
   873 => (x"c0",x"8c",x"78",x"c0"),
   874 => (x"c6",x"03",x"ac",x"b7"),
   875 => (x"a4",x"c0",x"c8",x"87"),
   876 => (x"c2",x"4c",x"c0",x"78"),
   877 => (x"bf",x"97",x"c7",x"dc"),
   878 => (x"02",x"99",x"d0",x"49"),
   879 => (x"1e",x"c0",x"87",x"d1"),
   880 => (x"49",x"cc",x"dc",x"c2"),
   881 => (x"c4",x"87",x"e4",x"eb"),
   882 => (x"4a",x"49",x"70",x"86"),
   883 => (x"c2",x"87",x"f6",x"c0"),
   884 => (x"c2",x"1e",x"d6",x"cf"),
   885 => (x"eb",x"49",x"cc",x"dc"),
   886 => (x"86",x"c4",x"87",x"d1"),
   887 => (x"ff",x"4a",x"49",x"70"),
   888 => (x"c5",x"c8",x"48",x"d0"),
   889 => (x"7b",x"d4",x"c1",x"78"),
   890 => (x"7b",x"bf",x"97",x"6e"),
   891 => (x"80",x"c1",x"48",x"6e"),
   892 => (x"66",x"c4",x"7e",x"70"),
   893 => (x"c8",x"88",x"c1",x"48"),
   894 => (x"98",x"70",x"58",x"a6"),
   895 => (x"87",x"e8",x"ff",x"05"),
   896 => (x"c4",x"48",x"d0",x"ff"),
   897 => (x"05",x"9a",x"72",x"78"),
   898 => (x"48",x"c0",x"87",x"c5"),
   899 => (x"c1",x"87",x"c2",x"c1"),
   900 => (x"cc",x"dc",x"c2",x"1e"),
   901 => (x"87",x"f9",x"e8",x"49"),
   902 => (x"9c",x"74",x"86",x"c4"),
   903 => (x"87",x"fc",x"fd",x"05"),
   904 => (x"06",x"ad",x"b7",x"c0"),
   905 => (x"dc",x"c2",x"87",x"d1"),
   906 => (x"78",x"c0",x"48",x"cc"),
   907 => (x"78",x"c0",x"80",x"d0"),
   908 => (x"dc",x"c2",x"80",x"f4"),
   909 => (x"c0",x"78",x"bf",x"d8"),
   910 => (x"fd",x"01",x"ad",x"b7"),
   911 => (x"d0",x"ff",x"87",x"d3"),
   912 => (x"c1",x"78",x"c5",x"48"),
   913 => (x"7b",x"c0",x"7b",x"d3"),
   914 => (x"48",x"c1",x"78",x"c4"),
   915 => (x"c0",x"87",x"c2",x"c0"),
   916 => (x"26",x"8e",x"f8",x"48"),
   917 => (x"26",x"4c",x"26",x"4d"),
   918 => (x"0e",x"4f",x"26",x"4b"),
   919 => (x"5d",x"5c",x"5b",x"5e"),
   920 => (x"4b",x"71",x"1e",x"0e"),
   921 => (x"ab",x"4d",x"4c",x"c0"),
   922 => (x"87",x"e8",x"c0",x"04"),
   923 => (x"1e",x"e5",x"f1",x"c0"),
   924 => (x"c4",x"02",x"9d",x"75"),
   925 => (x"c2",x"4a",x"c0",x"87"),
   926 => (x"72",x"4a",x"c1",x"87"),
   927 => (x"87",x"d0",x"ec",x"49"),
   928 => (x"7e",x"70",x"86",x"c4"),
   929 => (x"05",x"6e",x"84",x"c1"),
   930 => (x"4c",x"73",x"87",x"c2"),
   931 => (x"ac",x"73",x"85",x"c1"),
   932 => (x"87",x"d8",x"ff",x"06"),
   933 => (x"fe",x"26",x"48",x"6e"),
   934 => (x"71",x"1e",x"87",x"f9"),
   935 => (x"05",x"66",x"c4",x"4a"),
   936 => (x"49",x"72",x"87",x"c5"),
   937 => (x"26",x"87",x"de",x"f9"),
   938 => (x"5b",x"5e",x"0e",x"4f"),
   939 => (x"1e",x"0e",x"5d",x"5c"),
   940 => (x"de",x"49",x"4c",x"71"),
   941 => (x"f4",x"dc",x"c2",x"91"),
   942 => (x"97",x"85",x"71",x"4d"),
   943 => (x"dc",x"c1",x"02",x"6d"),
   944 => (x"e0",x"dc",x"c2",x"87"),
   945 => (x"82",x"74",x"4a",x"bf"),
   946 => (x"ce",x"fe",x"49",x"72"),
   947 => (x"6e",x"7e",x"70",x"87"),
   948 => (x"87",x"f2",x"c0",x"02"),
   949 => (x"4b",x"e8",x"dc",x"c2"),
   950 => (x"49",x"cb",x"4a",x"6e"),
   951 => (x"87",x"c8",x"c7",x"ff"),
   952 => (x"93",x"cb",x"4b",x"74"),
   953 => (x"83",x"f1",x"de",x"c1"),
   954 => (x"fc",x"c0",x"83",x"c4"),
   955 => (x"49",x"74",x"7b",x"e1"),
   956 => (x"87",x"de",x"c1",x"c1"),
   957 => (x"de",x"c1",x"7b",x"75"),
   958 => (x"49",x"bf",x"97",x"de"),
   959 => (x"e8",x"dc",x"c2",x"1e"),
   960 => (x"87",x"d6",x"fe",x"49"),
   961 => (x"49",x"74",x"86",x"c4"),
   962 => (x"87",x"c6",x"c1",x"c1"),
   963 => (x"c2",x"c1",x"49",x"c0"),
   964 => (x"dc",x"c2",x"87",x"e5"),
   965 => (x"78",x"c0",x"48",x"c8"),
   966 => (x"ea",x"de",x"49",x"c1"),
   967 => (x"f2",x"fc",x"26",x"87"),
   968 => (x"61",x"6f",x"4c",x"87"),
   969 => (x"67",x"6e",x"69",x"64"),
   970 => (x"00",x"2e",x"2e",x"2e"),
   971 => (x"5c",x"5b",x"5e",x"0e"),
   972 => (x"4a",x"4b",x"71",x"0e"),
   973 => (x"bf",x"e0",x"dc",x"c2"),
   974 => (x"fc",x"49",x"72",x"82"),
   975 => (x"4c",x"70",x"87",x"dd"),
   976 => (x"87",x"c4",x"02",x"9c"),
   977 => (x"87",x"d0",x"e8",x"49"),
   978 => (x"48",x"e0",x"dc",x"c2"),
   979 => (x"49",x"c1",x"78",x"c0"),
   980 => (x"fb",x"87",x"f4",x"dd"),
   981 => (x"c0",x"1e",x"87",x"ff"),
   982 => (x"da",x"c1",x"c1",x"49"),
   983 => (x"1e",x"4f",x"26",x"87"),
   984 => (x"cb",x"49",x"4a",x"71"),
   985 => (x"f1",x"de",x"c1",x"91"),
   986 => (x"11",x"81",x"c8",x"81"),
   987 => (x"cc",x"dc",x"c2",x"48"),
   988 => (x"e0",x"dc",x"c2",x"58"),
   989 => (x"c1",x"78",x"c0",x"48"),
   990 => (x"87",x"cb",x"dd",x"49"),
   991 => (x"71",x"1e",x"4f",x"26"),
   992 => (x"87",x"d2",x"02",x"99"),
   993 => (x"48",x"c6",x"e0",x"c1"),
   994 => (x"80",x"f7",x"50",x"c0"),
   995 => (x"40",x"df",x"fd",x"c0"),
   996 => (x"78",x"ea",x"de",x"c1"),
   997 => (x"e0",x"c1",x"87",x"ce"),
   998 => (x"de",x"c1",x"48",x"c2"),
   999 => (x"80",x"fc",x"78",x"e3"),
  1000 => (x"78",x"d6",x"fd",x"c0"),
  1001 => (x"5e",x"0e",x"4f",x"26"),
  1002 => (x"0e",x"5d",x"5c",x"5b"),
  1003 => (x"cf",x"c2",x"86",x"f4"),
  1004 => (x"4c",x"c0",x"4d",x"d6"),
  1005 => (x"c0",x"48",x"a6",x"c4"),
  1006 => (x"e0",x"dc",x"c2",x"78"),
  1007 => (x"a9",x"c0",x"49",x"bf"),
  1008 => (x"87",x"c1",x"c1",x"06"),
  1009 => (x"48",x"d6",x"cf",x"c2"),
  1010 => (x"f8",x"c0",x"02",x"98"),
  1011 => (x"e5",x"f1",x"c0",x"87"),
  1012 => (x"02",x"66",x"c8",x"1e"),
  1013 => (x"a6",x"c4",x"87",x"c7"),
  1014 => (x"c5",x"78",x"c0",x"48"),
  1015 => (x"48",x"a6",x"c4",x"87"),
  1016 => (x"66",x"c4",x"78",x"c1"),
  1017 => (x"87",x"e8",x"e6",x"49"),
  1018 => (x"4d",x"70",x"86",x"c4"),
  1019 => (x"66",x"c4",x"84",x"c1"),
  1020 => (x"c8",x"80",x"c1",x"48"),
  1021 => (x"dc",x"c2",x"58",x"a6"),
  1022 => (x"ac",x"49",x"bf",x"e0"),
  1023 => (x"75",x"87",x"c6",x"03"),
  1024 => (x"c8",x"ff",x"05",x"9d"),
  1025 => (x"75",x"4c",x"c0",x"87"),
  1026 => (x"e0",x"c3",x"02",x"9d"),
  1027 => (x"e5",x"f1",x"c0",x"87"),
  1028 => (x"02",x"66",x"c8",x"1e"),
  1029 => (x"a6",x"cc",x"87",x"c7"),
  1030 => (x"c5",x"78",x"c0",x"48"),
  1031 => (x"48",x"a6",x"cc",x"87"),
  1032 => (x"66",x"cc",x"78",x"c1"),
  1033 => (x"87",x"e8",x"e5",x"49"),
  1034 => (x"7e",x"70",x"86",x"c4"),
  1035 => (x"e9",x"c2",x"02",x"6e"),
  1036 => (x"cb",x"49",x"6e",x"87"),
  1037 => (x"49",x"69",x"97",x"81"),
  1038 => (x"c1",x"02",x"99",x"d0"),
  1039 => (x"fc",x"c0",x"87",x"d6"),
  1040 => (x"49",x"74",x"4a",x"ec"),
  1041 => (x"de",x"c1",x"91",x"cb"),
  1042 => (x"79",x"72",x"81",x"f1"),
  1043 => (x"ff",x"c3",x"81",x"c8"),
  1044 => (x"de",x"49",x"74",x"51"),
  1045 => (x"f4",x"dc",x"c2",x"91"),
  1046 => (x"c2",x"85",x"71",x"4d"),
  1047 => (x"c1",x"7d",x"97",x"c1"),
  1048 => (x"e0",x"c0",x"49",x"a5"),
  1049 => (x"e6",x"d7",x"c2",x"51"),
  1050 => (x"d2",x"02",x"bf",x"97"),
  1051 => (x"c2",x"84",x"c1",x"87"),
  1052 => (x"d7",x"c2",x"4b",x"a5"),
  1053 => (x"49",x"db",x"4a",x"e6"),
  1054 => (x"87",x"ec",x"c0",x"ff"),
  1055 => (x"cd",x"87",x"db",x"c1"),
  1056 => (x"51",x"c0",x"49",x"a5"),
  1057 => (x"a5",x"c2",x"84",x"c1"),
  1058 => (x"cb",x"4a",x"6e",x"4b"),
  1059 => (x"d7",x"c0",x"ff",x"49"),
  1060 => (x"87",x"c6",x"c1",x"87"),
  1061 => (x"4a",x"e9",x"fa",x"c0"),
  1062 => (x"91",x"cb",x"49",x"74"),
  1063 => (x"81",x"f1",x"de",x"c1"),
  1064 => (x"d7",x"c2",x"79",x"72"),
  1065 => (x"02",x"bf",x"97",x"e6"),
  1066 => (x"49",x"74",x"87",x"d8"),
  1067 => (x"84",x"c1",x"91",x"de"),
  1068 => (x"4b",x"f4",x"dc",x"c2"),
  1069 => (x"d7",x"c2",x"83",x"71"),
  1070 => (x"49",x"dd",x"4a",x"e6"),
  1071 => (x"87",x"e8",x"ff",x"fe"),
  1072 => (x"4b",x"74",x"87",x"d8"),
  1073 => (x"dc",x"c2",x"93",x"de"),
  1074 => (x"a3",x"cb",x"83",x"f4"),
  1075 => (x"c1",x"51",x"c0",x"49"),
  1076 => (x"4a",x"6e",x"73",x"84"),
  1077 => (x"ff",x"fe",x"49",x"cb"),
  1078 => (x"66",x"c4",x"87",x"ce"),
  1079 => (x"c8",x"80",x"c1",x"48"),
  1080 => (x"ac",x"c7",x"58",x"a6"),
  1081 => (x"87",x"c5",x"c0",x"03"),
  1082 => (x"e0",x"fc",x"05",x"6e"),
  1083 => (x"f4",x"48",x"74",x"87"),
  1084 => (x"87",x"df",x"f5",x"8e"),
  1085 => (x"71",x"1e",x"73",x"1e"),
  1086 => (x"91",x"cb",x"49",x"4b"),
  1087 => (x"81",x"f1",x"de",x"c1"),
  1088 => (x"c1",x"4a",x"a1",x"c8"),
  1089 => (x"12",x"48",x"dd",x"de"),
  1090 => (x"4a",x"a1",x"c9",x"50"),
  1091 => (x"48",x"c4",x"f4",x"c0"),
  1092 => (x"81",x"ca",x"50",x"12"),
  1093 => (x"48",x"de",x"de",x"c1"),
  1094 => (x"de",x"c1",x"50",x"11"),
  1095 => (x"49",x"bf",x"97",x"de"),
  1096 => (x"f5",x"49",x"c0",x"1e"),
  1097 => (x"dc",x"c2",x"87",x"f4"),
  1098 => (x"78",x"de",x"48",x"c8"),
  1099 => (x"d6",x"d6",x"49",x"c1"),
  1100 => (x"e2",x"f4",x"26",x"87"),
  1101 => (x"5b",x"5e",x"0e",x"87"),
  1102 => (x"f4",x"0e",x"5d",x"5c"),
  1103 => (x"49",x"4d",x"71",x"86"),
  1104 => (x"de",x"c1",x"91",x"cb"),
  1105 => (x"a1",x"c8",x"81",x"f1"),
  1106 => (x"7e",x"a1",x"ca",x"4a"),
  1107 => (x"c2",x"48",x"a6",x"c4"),
  1108 => (x"78",x"bf",x"d0",x"e0"),
  1109 => (x"4b",x"bf",x"97",x"6e"),
  1110 => (x"73",x"48",x"66",x"c4"),
  1111 => (x"4c",x"4b",x"70",x"28"),
  1112 => (x"a6",x"cc",x"48",x"12"),
  1113 => (x"c1",x"9c",x"70",x"58"),
  1114 => (x"97",x"81",x"c9",x"84"),
  1115 => (x"ac",x"b7",x"49",x"69"),
  1116 => (x"c0",x"87",x"c2",x"04"),
  1117 => (x"bf",x"97",x"6e",x"4c"),
  1118 => (x"49",x"66",x"c8",x"4a"),
  1119 => (x"b9",x"ff",x"31",x"72"),
  1120 => (x"74",x"99",x"66",x"c4"),
  1121 => (x"70",x"30",x"72",x"48"),
  1122 => (x"b0",x"71",x"48",x"4a"),
  1123 => (x"58",x"d4",x"e0",x"c2"),
  1124 => (x"87",x"fe",x"e4",x"c0"),
  1125 => (x"ee",x"d4",x"49",x"c0"),
  1126 => (x"c0",x"49",x"75",x"87"),
  1127 => (x"f4",x"87",x"f3",x"f6"),
  1128 => (x"87",x"ef",x"f2",x"8e"),
  1129 => (x"71",x"1e",x"73",x"1e"),
  1130 => (x"c8",x"fe",x"49",x"4b"),
  1131 => (x"fe",x"49",x"73",x"87"),
  1132 => (x"e2",x"f2",x"87",x"c3"),
  1133 => (x"1e",x"73",x"1e",x"87"),
  1134 => (x"a3",x"c6",x"4b",x"71"),
  1135 => (x"e3",x"c0",x"02",x"4a"),
  1136 => (x"02",x"8a",x"c1",x"87"),
  1137 => (x"02",x"8a",x"87",x"d6"),
  1138 => (x"8a",x"87",x"e8",x"c1"),
  1139 => (x"87",x"ca",x"c1",x"02"),
  1140 => (x"ef",x"c0",x"02",x"8a"),
  1141 => (x"d9",x"02",x"8a",x"87"),
  1142 => (x"87",x"e9",x"c1",x"87"),
  1143 => (x"fe",x"f5",x"49",x"c7"),
  1144 => (x"87",x"ec",x"c1",x"87"),
  1145 => (x"48",x"c8",x"dc",x"c2"),
  1146 => (x"49",x"c1",x"78",x"df"),
  1147 => (x"c1",x"87",x"d8",x"d3"),
  1148 => (x"dc",x"c2",x"87",x"de"),
  1149 => (x"c1",x"02",x"bf",x"e0"),
  1150 => (x"c1",x"48",x"87",x"cb"),
  1151 => (x"e4",x"dc",x"c2",x"88"),
  1152 => (x"87",x"c1",x"c1",x"58"),
  1153 => (x"bf",x"e4",x"dc",x"c2"),
  1154 => (x"87",x"f9",x"c0",x"02"),
  1155 => (x"bf",x"e0",x"dc",x"c2"),
  1156 => (x"c2",x"80",x"c1",x"48"),
  1157 => (x"c0",x"58",x"e4",x"dc"),
  1158 => (x"dc",x"c2",x"87",x"eb"),
  1159 => (x"c6",x"49",x"bf",x"e0"),
  1160 => (x"e4",x"dc",x"c2",x"89"),
  1161 => (x"a9",x"b7",x"c0",x"59"),
  1162 => (x"c2",x"87",x"da",x"03"),
  1163 => (x"c0",x"48",x"e0",x"dc"),
  1164 => (x"c2",x"87",x"d2",x"78"),
  1165 => (x"02",x"bf",x"e4",x"dc"),
  1166 => (x"dc",x"c2",x"87",x"cb"),
  1167 => (x"c6",x"48",x"bf",x"e0"),
  1168 => (x"e4",x"dc",x"c2",x"80"),
  1169 => (x"d1",x"49",x"c0",x"58"),
  1170 => (x"49",x"73",x"87",x"fd"),
  1171 => (x"87",x"c2",x"f4",x"c0"),
  1172 => (x"0e",x"87",x"c4",x"f0"),
  1173 => (x"5d",x"5c",x"5b",x"5e"),
  1174 => (x"86",x"d0",x"ff",x"0e"),
  1175 => (x"c8",x"59",x"a6",x"dc"),
  1176 => (x"78",x"c0",x"48",x"a6"),
  1177 => (x"c4",x"c1",x"80",x"c4"),
  1178 => (x"80",x"c4",x"78",x"66"),
  1179 => (x"80",x"c4",x"78",x"c1"),
  1180 => (x"dc",x"c2",x"78",x"c1"),
  1181 => (x"78",x"c1",x"48",x"e4"),
  1182 => (x"bf",x"c8",x"dc",x"c2"),
  1183 => (x"05",x"a8",x"de",x"48"),
  1184 => (x"e1",x"f4",x"87",x"cb"),
  1185 => (x"cc",x"49",x"70",x"87"),
  1186 => (x"f9",x"cf",x"59",x"a6"),
  1187 => (x"87",x"c4",x"e4",x"87"),
  1188 => (x"e3",x"87",x"e6",x"e4"),
  1189 => (x"4c",x"70",x"87",x"f3"),
  1190 => (x"02",x"ac",x"fb",x"c0"),
  1191 => (x"d8",x"87",x"fb",x"c1"),
  1192 => (x"ed",x"c1",x"05",x"66"),
  1193 => (x"66",x"c0",x"c1",x"87"),
  1194 => (x"6a",x"82",x"c4",x"4a"),
  1195 => (x"c1",x"1e",x"72",x"7e"),
  1196 => (x"c4",x"48",x"fb",x"da"),
  1197 => (x"a1",x"c8",x"49",x"66"),
  1198 => (x"71",x"41",x"20",x"4a"),
  1199 => (x"87",x"f9",x"05",x"aa"),
  1200 => (x"4a",x"26",x"51",x"10"),
  1201 => (x"48",x"66",x"c0",x"c1"),
  1202 => (x"78",x"f4",x"c3",x"c1"),
  1203 => (x"81",x"c7",x"49",x"6a"),
  1204 => (x"c0",x"c1",x"51",x"74"),
  1205 => (x"81",x"c8",x"49",x"66"),
  1206 => (x"c0",x"c1",x"51",x"c1"),
  1207 => (x"81",x"c9",x"49",x"66"),
  1208 => (x"c0",x"c1",x"51",x"c0"),
  1209 => (x"81",x"ca",x"49",x"66"),
  1210 => (x"1e",x"c1",x"51",x"c0"),
  1211 => (x"49",x"6a",x"1e",x"d8"),
  1212 => (x"d8",x"e3",x"81",x"c8"),
  1213 => (x"c1",x"86",x"c8",x"87"),
  1214 => (x"c0",x"48",x"66",x"c4"),
  1215 => (x"87",x"c7",x"01",x"a8"),
  1216 => (x"c1",x"48",x"a6",x"c8"),
  1217 => (x"c1",x"87",x"ce",x"78"),
  1218 => (x"c1",x"48",x"66",x"c4"),
  1219 => (x"58",x"a6",x"d0",x"88"),
  1220 => (x"e4",x"e2",x"87",x"c3"),
  1221 => (x"48",x"a6",x"d0",x"87"),
  1222 => (x"9c",x"74",x"78",x"c2"),
  1223 => (x"87",x"e2",x"cd",x"02"),
  1224 => (x"c1",x"48",x"66",x"c8"),
  1225 => (x"03",x"a8",x"66",x"c8"),
  1226 => (x"dc",x"87",x"d7",x"cd"),
  1227 => (x"78",x"c0",x"48",x"a6"),
  1228 => (x"78",x"c0",x"80",x"e8"),
  1229 => (x"70",x"87",x"d2",x"e1"),
  1230 => (x"ac",x"d0",x"c1",x"4c"),
  1231 => (x"87",x"d7",x"c2",x"05"),
  1232 => (x"e3",x"7e",x"66",x"c4"),
  1233 => (x"49",x"70",x"87",x"f6"),
  1234 => (x"e0",x"59",x"a6",x"c8"),
  1235 => (x"4c",x"70",x"87",x"fb"),
  1236 => (x"05",x"ac",x"ec",x"c0"),
  1237 => (x"c8",x"87",x"eb",x"c1"),
  1238 => (x"91",x"cb",x"49",x"66"),
  1239 => (x"81",x"66",x"c0",x"c1"),
  1240 => (x"6a",x"4a",x"a1",x"c4"),
  1241 => (x"4a",x"a1",x"c8",x"4d"),
  1242 => (x"c0",x"52",x"66",x"c4"),
  1243 => (x"e0",x"79",x"df",x"fd"),
  1244 => (x"4c",x"70",x"87",x"d7"),
  1245 => (x"87",x"d8",x"02",x"9c"),
  1246 => (x"02",x"ac",x"fb",x"c0"),
  1247 => (x"55",x"74",x"87",x"d2"),
  1248 => (x"70",x"87",x"c6",x"e0"),
  1249 => (x"c7",x"02",x"9c",x"4c"),
  1250 => (x"ac",x"fb",x"c0",x"87"),
  1251 => (x"87",x"ee",x"ff",x"05"),
  1252 => (x"c2",x"55",x"e0",x"c0"),
  1253 => (x"97",x"c0",x"55",x"c1"),
  1254 => (x"49",x"66",x"d8",x"7d"),
  1255 => (x"db",x"05",x"a9",x"6e"),
  1256 => (x"48",x"66",x"c8",x"87"),
  1257 => (x"04",x"a8",x"66",x"cc"),
  1258 => (x"66",x"c8",x"87",x"ca"),
  1259 => (x"cc",x"80",x"c1",x"48"),
  1260 => (x"87",x"c8",x"58",x"a6"),
  1261 => (x"c1",x"48",x"66",x"cc"),
  1262 => (x"58",x"a6",x"d0",x"88"),
  1263 => (x"87",x"c9",x"df",x"ff"),
  1264 => (x"d0",x"c1",x"4c",x"70"),
  1265 => (x"87",x"c8",x"05",x"ac"),
  1266 => (x"c1",x"48",x"66",x"d4"),
  1267 => (x"58",x"a6",x"d8",x"80"),
  1268 => (x"02",x"ac",x"d0",x"c1"),
  1269 => (x"c0",x"87",x"e9",x"fd"),
  1270 => (x"d8",x"48",x"a6",x"e0"),
  1271 => (x"66",x"c4",x"78",x"66"),
  1272 => (x"66",x"e0",x"c0",x"48"),
  1273 => (x"eb",x"c9",x"05",x"a8"),
  1274 => (x"a6",x"e4",x"c0",x"87"),
  1275 => (x"74",x"78",x"c0",x"48"),
  1276 => (x"88",x"fb",x"c0",x"48"),
  1277 => (x"02",x"6e",x"7e",x"70"),
  1278 => (x"6e",x"87",x"ee",x"c9"),
  1279 => (x"70",x"88",x"cb",x"48"),
  1280 => (x"c1",x"02",x"6e",x"7e"),
  1281 => (x"48",x"6e",x"87",x"cd"),
  1282 => (x"7e",x"70",x"88",x"c9"),
  1283 => (x"c1",x"c4",x"02",x"6e"),
  1284 => (x"c4",x"48",x"6e",x"87"),
  1285 => (x"6e",x"7e",x"70",x"88"),
  1286 => (x"6e",x"87",x"ce",x"02"),
  1287 => (x"70",x"88",x"c1",x"48"),
  1288 => (x"c3",x"02",x"6e",x"7e"),
  1289 => (x"e2",x"c8",x"87",x"ec"),
  1290 => (x"48",x"a6",x"dc",x"87"),
  1291 => (x"ff",x"78",x"f0",x"c0"),
  1292 => (x"70",x"87",x"d6",x"dd"),
  1293 => (x"ac",x"ec",x"c0",x"4c"),
  1294 => (x"87",x"c4",x"c0",x"02"),
  1295 => (x"5c",x"a6",x"e0",x"c0"),
  1296 => (x"02",x"ac",x"ec",x"c0"),
  1297 => (x"dc",x"ff",x"87",x"cd"),
  1298 => (x"4c",x"70",x"87",x"ff"),
  1299 => (x"05",x"ac",x"ec",x"c0"),
  1300 => (x"c0",x"87",x"f3",x"ff"),
  1301 => (x"c0",x"02",x"ac",x"ec"),
  1302 => (x"dc",x"ff",x"87",x"c4"),
  1303 => (x"1e",x"c0",x"87",x"eb"),
  1304 => (x"66",x"d0",x"1e",x"ca"),
  1305 => (x"c1",x"91",x"cb",x"49"),
  1306 => (x"71",x"48",x"66",x"c8"),
  1307 => (x"58",x"a6",x"cc",x"80"),
  1308 => (x"c4",x"48",x"66",x"c8"),
  1309 => (x"58",x"a6",x"d0",x"80"),
  1310 => (x"49",x"bf",x"66",x"cc"),
  1311 => (x"87",x"cd",x"dd",x"ff"),
  1312 => (x"1e",x"de",x"1e",x"c1"),
  1313 => (x"49",x"bf",x"66",x"d4"),
  1314 => (x"87",x"c1",x"dd",x"ff"),
  1315 => (x"49",x"70",x"86",x"d0"),
  1316 => (x"c0",x"89",x"09",x"c0"),
  1317 => (x"c0",x"59",x"a6",x"ec"),
  1318 => (x"c0",x"48",x"66",x"e8"),
  1319 => (x"ee",x"c0",x"06",x"a8"),
  1320 => (x"66",x"e8",x"c0",x"87"),
  1321 => (x"03",x"a8",x"dd",x"48"),
  1322 => (x"c4",x"87",x"e4",x"c0"),
  1323 => (x"c0",x"49",x"bf",x"66"),
  1324 => (x"c0",x"81",x"66",x"e8"),
  1325 => (x"e8",x"c0",x"51",x"e0"),
  1326 => (x"81",x"c1",x"49",x"66"),
  1327 => (x"81",x"bf",x"66",x"c4"),
  1328 => (x"c0",x"51",x"c1",x"c2"),
  1329 => (x"c2",x"49",x"66",x"e8"),
  1330 => (x"bf",x"66",x"c4",x"81"),
  1331 => (x"6e",x"51",x"c0",x"81"),
  1332 => (x"f4",x"c3",x"c1",x"48"),
  1333 => (x"c8",x"49",x"6e",x"78"),
  1334 => (x"51",x"66",x"d0",x"81"),
  1335 => (x"81",x"c9",x"49",x"6e"),
  1336 => (x"6e",x"51",x"66",x"d4"),
  1337 => (x"dc",x"81",x"ca",x"49"),
  1338 => (x"66",x"d0",x"51",x"66"),
  1339 => (x"d4",x"80",x"c1",x"48"),
  1340 => (x"66",x"c8",x"58",x"a6"),
  1341 => (x"a8",x"66",x"cc",x"48"),
  1342 => (x"87",x"cb",x"c0",x"04"),
  1343 => (x"c1",x"48",x"66",x"c8"),
  1344 => (x"58",x"a6",x"cc",x"80"),
  1345 => (x"cc",x"87",x"e2",x"c5"),
  1346 => (x"88",x"c1",x"48",x"66"),
  1347 => (x"c5",x"58",x"a6",x"d0"),
  1348 => (x"dc",x"ff",x"87",x"d7"),
  1349 => (x"49",x"70",x"87",x"e6"),
  1350 => (x"59",x"a6",x"ec",x"c0"),
  1351 => (x"87",x"dc",x"dc",x"ff"),
  1352 => (x"e0",x"c0",x"49",x"70"),
  1353 => (x"66",x"dc",x"59",x"a6"),
  1354 => (x"a8",x"ec",x"c0",x"48"),
  1355 => (x"87",x"ca",x"c0",x"05"),
  1356 => (x"c0",x"48",x"a6",x"dc"),
  1357 => (x"c0",x"78",x"66",x"e8"),
  1358 => (x"d9",x"ff",x"87",x"c4"),
  1359 => (x"66",x"c8",x"87",x"cb"),
  1360 => (x"c1",x"91",x"cb",x"49"),
  1361 => (x"71",x"48",x"66",x"c0"),
  1362 => (x"6e",x"7e",x"70",x"80"),
  1363 => (x"6e",x"82",x"c8",x"4a"),
  1364 => (x"c0",x"81",x"ca",x"49"),
  1365 => (x"dc",x"51",x"66",x"e8"),
  1366 => (x"81",x"c1",x"49",x"66"),
  1367 => (x"89",x"66",x"e8",x"c0"),
  1368 => (x"30",x"71",x"48",x"c1"),
  1369 => (x"89",x"c1",x"49",x"70"),
  1370 => (x"c2",x"7a",x"97",x"71"),
  1371 => (x"49",x"bf",x"d0",x"e0"),
  1372 => (x"29",x"66",x"e8",x"c0"),
  1373 => (x"48",x"4a",x"6a",x"97"),
  1374 => (x"f0",x"c0",x"98",x"71"),
  1375 => (x"49",x"6e",x"58",x"a6"),
  1376 => (x"4d",x"69",x"81",x"c4"),
  1377 => (x"48",x"66",x"e0",x"c0"),
  1378 => (x"02",x"a8",x"66",x"c4"),
  1379 => (x"c4",x"87",x"c8",x"c0"),
  1380 => (x"78",x"c0",x"48",x"a6"),
  1381 => (x"c4",x"87",x"c5",x"c0"),
  1382 => (x"78",x"c1",x"48",x"a6"),
  1383 => (x"c0",x"1e",x"66",x"c4"),
  1384 => (x"49",x"75",x"1e",x"e0"),
  1385 => (x"87",x"e5",x"d8",x"ff"),
  1386 => (x"4c",x"70",x"86",x"c8"),
  1387 => (x"06",x"ac",x"b7",x"c0"),
  1388 => (x"74",x"87",x"d4",x"c1"),
  1389 => (x"49",x"e0",x"c0",x"85"),
  1390 => (x"4b",x"75",x"89",x"74"),
  1391 => (x"4a",x"c4",x"db",x"c1"),
  1392 => (x"e3",x"eb",x"fe",x"71"),
  1393 => (x"c0",x"85",x"c2",x"87"),
  1394 => (x"c1",x"48",x"66",x"e4"),
  1395 => (x"a6",x"e8",x"c0",x"80"),
  1396 => (x"66",x"ec",x"c0",x"58"),
  1397 => (x"70",x"81",x"c1",x"49"),
  1398 => (x"c8",x"c0",x"02",x"a9"),
  1399 => (x"48",x"a6",x"c4",x"87"),
  1400 => (x"c5",x"c0",x"78",x"c0"),
  1401 => (x"48",x"a6",x"c4",x"87"),
  1402 => (x"66",x"c4",x"78",x"c1"),
  1403 => (x"49",x"a4",x"c2",x"1e"),
  1404 => (x"71",x"48",x"e0",x"c0"),
  1405 => (x"1e",x"49",x"70",x"88"),
  1406 => (x"d7",x"ff",x"49",x"75"),
  1407 => (x"86",x"c8",x"87",x"cf"),
  1408 => (x"01",x"a8",x"b7",x"c0"),
  1409 => (x"c0",x"87",x"c0",x"ff"),
  1410 => (x"c0",x"02",x"66",x"e4"),
  1411 => (x"49",x"6e",x"87",x"d1"),
  1412 => (x"e4",x"c0",x"81",x"c9"),
  1413 => (x"48",x"6e",x"51",x"66"),
  1414 => (x"78",x"f5",x"c4",x"c1"),
  1415 => (x"6e",x"87",x"cc",x"c0"),
  1416 => (x"c2",x"81",x"c9",x"49"),
  1417 => (x"c1",x"48",x"6e",x"51"),
  1418 => (x"c8",x"78",x"e4",x"c6"),
  1419 => (x"66",x"cc",x"48",x"66"),
  1420 => (x"cb",x"c0",x"04",x"a8"),
  1421 => (x"48",x"66",x"c8",x"87"),
  1422 => (x"a6",x"cc",x"80",x"c1"),
  1423 => (x"87",x"e9",x"c0",x"58"),
  1424 => (x"c1",x"48",x"66",x"cc"),
  1425 => (x"58",x"a6",x"d0",x"88"),
  1426 => (x"ff",x"87",x"de",x"c0"),
  1427 => (x"70",x"87",x"ea",x"d5"),
  1428 => (x"87",x"d5",x"c0",x"4c"),
  1429 => (x"05",x"ac",x"c6",x"c1"),
  1430 => (x"d0",x"87",x"c8",x"c0"),
  1431 => (x"80",x"c1",x"48",x"66"),
  1432 => (x"ff",x"58",x"a6",x"d4"),
  1433 => (x"70",x"87",x"d2",x"d5"),
  1434 => (x"48",x"66",x"d4",x"4c"),
  1435 => (x"a6",x"d8",x"80",x"c1"),
  1436 => (x"02",x"9c",x"74",x"58"),
  1437 => (x"c8",x"87",x"cb",x"c0"),
  1438 => (x"c8",x"c1",x"48",x"66"),
  1439 => (x"f2",x"04",x"a8",x"66"),
  1440 => (x"d4",x"ff",x"87",x"e9"),
  1441 => (x"66",x"c8",x"87",x"ea"),
  1442 => (x"03",x"a8",x"c7",x"48"),
  1443 => (x"c2",x"87",x"e5",x"c0"),
  1444 => (x"c0",x"48",x"e4",x"dc"),
  1445 => (x"49",x"66",x"c8",x"78"),
  1446 => (x"c0",x"c1",x"91",x"cb"),
  1447 => (x"a1",x"c4",x"81",x"66"),
  1448 => (x"c0",x"4a",x"6a",x"4a"),
  1449 => (x"66",x"c8",x"79",x"52"),
  1450 => (x"cc",x"80",x"c1",x"48"),
  1451 => (x"a8",x"c7",x"58",x"a6"),
  1452 => (x"87",x"db",x"ff",x"04"),
  1453 => (x"ff",x"8e",x"d0",x"ff"),
  1454 => (x"4c",x"87",x"d8",x"de"),
  1455 => (x"20",x"64",x"61",x"6f"),
  1456 => (x"00",x"20",x"2e",x"2a"),
  1457 => (x"1e",x"00",x"20",x"3a"),
  1458 => (x"4b",x"71",x"1e",x"73"),
  1459 => (x"87",x"c6",x"02",x"9b"),
  1460 => (x"48",x"e0",x"dc",x"c2"),
  1461 => (x"1e",x"c7",x"78",x"c0"),
  1462 => (x"bf",x"e0",x"dc",x"c2"),
  1463 => (x"de",x"c1",x"1e",x"49"),
  1464 => (x"dc",x"c2",x"1e",x"f1"),
  1465 => (x"ed",x"49",x"bf",x"c8"),
  1466 => (x"86",x"cc",x"87",x"e9"),
  1467 => (x"bf",x"c8",x"dc",x"c2"),
  1468 => (x"87",x"ca",x"e2",x"49"),
  1469 => (x"c8",x"02",x"9b",x"73"),
  1470 => (x"f1",x"de",x"c1",x"87"),
  1471 => (x"e3",x"e2",x"c0",x"49"),
  1472 => (x"d2",x"dd",x"ff",x"87"),
  1473 => (x"de",x"c1",x"1e",x"87"),
  1474 => (x"50",x"c0",x"48",x"dd"),
  1475 => (x"bf",x"d4",x"e0",x"c1"),
  1476 => (x"f0",x"d7",x"ff",x"49"),
  1477 => (x"26",x"48",x"c0",x"87"),
  1478 => (x"de",x"c7",x"1e",x"4f"),
  1479 => (x"fe",x"49",x"c1",x"87"),
  1480 => (x"ee",x"fe",x"87",x"e5"),
  1481 => (x"98",x"70",x"87",x"c3"),
  1482 => (x"fe",x"87",x"cd",x"02"),
  1483 => (x"70",x"87",x"dc",x"f5"),
  1484 => (x"87",x"c4",x"02",x"98"),
  1485 => (x"87",x"c2",x"4a",x"c1"),
  1486 => (x"9a",x"72",x"4a",x"c0"),
  1487 => (x"c0",x"87",x"ce",x"05"),
  1488 => (x"f4",x"dd",x"c1",x"1e"),
  1489 => (x"e0",x"ef",x"c0",x"49"),
  1490 => (x"fe",x"86",x"c4",x"87"),
  1491 => (x"e0",x"dc",x"c2",x"87"),
  1492 => (x"c2",x"78",x"c0",x"48"),
  1493 => (x"c0",x"48",x"c8",x"dc"),
  1494 => (x"dd",x"c1",x"1e",x"78"),
  1495 => (x"ef",x"c0",x"49",x"ff"),
  1496 => (x"1e",x"c0",x"87",x"c7"),
  1497 => (x"70",x"87",x"de",x"fe"),
  1498 => (x"fc",x"ee",x"c0",x"49"),
  1499 => (x"87",x"ca",x"c3",x"87"),
  1500 => (x"4f",x"26",x"8e",x"f8"),
  1501 => (x"66",x"20",x"44",x"53"),
  1502 => (x"65",x"6c",x"69",x"61"),
  1503 => (x"42",x"00",x"2e",x"64"),
  1504 => (x"69",x"74",x"6f",x"6f"),
  1505 => (x"2e",x"2e",x"67",x"6e"),
  1506 => (x"c0",x"1e",x"00",x"2e"),
  1507 => (x"fa",x"87",x"d2",x"e2"),
  1508 => (x"1e",x"4f",x"26",x"87"),
  1509 => (x"f1",x"87",x"c2",x"fe"),
  1510 => (x"26",x"48",x"c0",x"87"),
  1511 => (x"01",x"00",x"00",x"4f"),
  1512 => (x"80",x"00",x"00",x"00"),
  1513 => (x"69",x"78",x"45",x"20"),
  1514 => (x"20",x"80",x"00",x"74"),
  1515 => (x"6b",x"63",x"61",x"42"),
  1516 => (x"00",x"0e",x"a9",x"00"),
  1517 => (x"00",x"27",x"34",x"00"),
  1518 => (x"00",x"00",x"00",x"00"),
  1519 => (x"00",x"00",x"0e",x"a9"),
  1520 => (x"00",x"00",x"27",x"52"),
  1521 => (x"a9",x"00",x"00",x"00"),
  1522 => (x"70",x"00",x"00",x"0e"),
  1523 => (x"00",x"00",x"00",x"27"),
  1524 => (x"0e",x"a9",x"00",x"00"),
  1525 => (x"27",x"8e",x"00",x"00"),
  1526 => (x"00",x"00",x"00",x"00"),
  1527 => (x"00",x"0e",x"a9",x"00"),
  1528 => (x"00",x"27",x"ac",x"00"),
  1529 => (x"00",x"00",x"00",x"00"),
  1530 => (x"00",x"00",x"0e",x"a9"),
  1531 => (x"00",x"00",x"27",x"ca"),
  1532 => (x"a9",x"00",x"00",x"00"),
  1533 => (x"e8",x"00",x"00",x"0e"),
  1534 => (x"00",x"00",x"00",x"27"),
  1535 => (x"0f",x"5f",x"00",x"00"),
  1536 => (x"00",x"00",x"00",x"00"),
  1537 => (x"00",x"00",x"00",x"00"),
  1538 => (x"00",x"11",x"b5",x"00"),
  1539 => (x"00",x"00",x"00",x"00"),
  1540 => (x"00",x"00",x"00",x"00"),
  1541 => (x"00",x"00",x"18",x"18"),
  1542 => (x"54",x"4f",x"4f",x"42"),
  1543 => (x"20",x"20",x"20",x"20"),
  1544 => (x"00",x"4d",x"4f",x"52"),
  1545 => (x"48",x"f0",x"fe",x"1e"),
  1546 => (x"09",x"cd",x"78",x"c0"),
  1547 => (x"4f",x"26",x"09",x"79"),
  1548 => (x"f0",x"fe",x"1e",x"1e"),
  1549 => (x"26",x"48",x"7e",x"bf"),
  1550 => (x"fe",x"1e",x"4f",x"26"),
  1551 => (x"78",x"c1",x"48",x"f0"),
  1552 => (x"fe",x"1e",x"4f",x"26"),
  1553 => (x"78",x"c0",x"48",x"f0"),
  1554 => (x"71",x"1e",x"4f",x"26"),
  1555 => (x"52",x"52",x"c0",x"4a"),
  1556 => (x"5e",x"0e",x"4f",x"26"),
  1557 => (x"0e",x"5d",x"5c",x"5b"),
  1558 => (x"4d",x"71",x"86",x"f4"),
  1559 => (x"c1",x"7e",x"6d",x"97"),
  1560 => (x"6c",x"97",x"4c",x"a5"),
  1561 => (x"58",x"a6",x"c8",x"48"),
  1562 => (x"66",x"c4",x"48",x"6e"),
  1563 => (x"87",x"c5",x"05",x"a8"),
  1564 => (x"e6",x"c0",x"48",x"ff"),
  1565 => (x"87",x"ca",x"ff",x"87"),
  1566 => (x"97",x"49",x"a5",x"c2"),
  1567 => (x"a3",x"71",x"4b",x"6c"),
  1568 => (x"4b",x"6b",x"97",x"4b"),
  1569 => (x"6e",x"7e",x"6c",x"97"),
  1570 => (x"c8",x"80",x"c1",x"48"),
  1571 => (x"98",x"c7",x"58",x"a6"),
  1572 => (x"70",x"58",x"a6",x"cc"),
  1573 => (x"e1",x"fe",x"7c",x"97"),
  1574 => (x"f4",x"48",x"73",x"87"),
  1575 => (x"26",x"4d",x"26",x"8e"),
  1576 => (x"26",x"4b",x"26",x"4c"),
  1577 => (x"5b",x"5e",x"0e",x"4f"),
  1578 => (x"86",x"f4",x"0e",x"5c"),
  1579 => (x"66",x"d8",x"4c",x"71"),
  1580 => (x"9a",x"ff",x"c3",x"4a"),
  1581 => (x"97",x"4b",x"a4",x"c2"),
  1582 => (x"a1",x"73",x"49",x"6c"),
  1583 => (x"97",x"51",x"72",x"49"),
  1584 => (x"48",x"6e",x"7e",x"6c"),
  1585 => (x"a6",x"c8",x"80",x"c1"),
  1586 => (x"cc",x"98",x"c7",x"58"),
  1587 => (x"54",x"70",x"58",x"a6"),
  1588 => (x"ca",x"ff",x"8e",x"f4"),
  1589 => (x"fd",x"1e",x"1e",x"87"),
  1590 => (x"bf",x"e0",x"87",x"e8"),
  1591 => (x"e0",x"c0",x"49",x"4a"),
  1592 => (x"cb",x"02",x"99",x"c0"),
  1593 => (x"c2",x"1e",x"72",x"87"),
  1594 => (x"fe",x"49",x"c6",x"e0"),
  1595 => (x"86",x"c4",x"87",x"f7"),
  1596 => (x"70",x"87",x"fd",x"fc"),
  1597 => (x"87",x"c2",x"fd",x"7e"),
  1598 => (x"1e",x"4f",x"26",x"26"),
  1599 => (x"49",x"c6",x"e0",x"c2"),
  1600 => (x"c1",x"87",x"c7",x"fd"),
  1601 => (x"fc",x"49",x"d5",x"e3"),
  1602 => (x"ee",x"c3",x"87",x"da"),
  1603 => (x"0e",x"4f",x"26",x"87"),
  1604 => (x"5d",x"5c",x"5b",x"5e"),
  1605 => (x"c2",x"4d",x"71",x"0e"),
  1606 => (x"fc",x"49",x"c6",x"e0"),
  1607 => (x"4b",x"70",x"87",x"f4"),
  1608 => (x"04",x"ab",x"b7",x"c0"),
  1609 => (x"c3",x"87",x"c2",x"c3"),
  1610 => (x"c9",x"05",x"ab",x"f0"),
  1611 => (x"f3",x"e7",x"c1",x"87"),
  1612 => (x"c2",x"78",x"c1",x"48"),
  1613 => (x"e0",x"c3",x"87",x"e3"),
  1614 => (x"87",x"c9",x"05",x"ab"),
  1615 => (x"48",x"f7",x"e7",x"c1"),
  1616 => (x"d4",x"c2",x"78",x"c1"),
  1617 => (x"f7",x"e7",x"c1",x"87"),
  1618 => (x"87",x"c6",x"02",x"bf"),
  1619 => (x"4c",x"a3",x"c0",x"c2"),
  1620 => (x"4c",x"73",x"87",x"c2"),
  1621 => (x"bf",x"f3",x"e7",x"c1"),
  1622 => (x"87",x"e0",x"c0",x"02"),
  1623 => (x"b7",x"c4",x"49",x"74"),
  1624 => (x"e9",x"c1",x"91",x"29"),
  1625 => (x"4a",x"74",x"81",x"ca"),
  1626 => (x"92",x"c2",x"9a",x"cf"),
  1627 => (x"30",x"72",x"48",x"c1"),
  1628 => (x"ba",x"ff",x"4a",x"70"),
  1629 => (x"98",x"69",x"48",x"72"),
  1630 => (x"87",x"db",x"79",x"70"),
  1631 => (x"b7",x"c4",x"49",x"74"),
  1632 => (x"e9",x"c1",x"91",x"29"),
  1633 => (x"4a",x"74",x"81",x"ca"),
  1634 => (x"92",x"c2",x"9a",x"cf"),
  1635 => (x"30",x"72",x"48",x"c3"),
  1636 => (x"69",x"48",x"4a",x"70"),
  1637 => (x"75",x"79",x"70",x"b0"),
  1638 => (x"f0",x"c0",x"05",x"9d"),
  1639 => (x"48",x"d0",x"ff",x"87"),
  1640 => (x"ff",x"78",x"e1",x"c8"),
  1641 => (x"78",x"c5",x"48",x"d4"),
  1642 => (x"bf",x"f7",x"e7",x"c1"),
  1643 => (x"c3",x"87",x"c3",x"02"),
  1644 => (x"e7",x"c1",x"78",x"e0"),
  1645 => (x"c6",x"02",x"bf",x"f3"),
  1646 => (x"48",x"d4",x"ff",x"87"),
  1647 => (x"ff",x"78",x"f0",x"c3"),
  1648 => (x"78",x"73",x"48",x"d4"),
  1649 => (x"c8",x"48",x"d0",x"ff"),
  1650 => (x"e0",x"c0",x"78",x"e1"),
  1651 => (x"f7",x"e7",x"c1",x"78"),
  1652 => (x"c1",x"78",x"c0",x"48"),
  1653 => (x"c0",x"48",x"f3",x"e7"),
  1654 => (x"c6",x"e0",x"c2",x"78"),
  1655 => (x"87",x"f2",x"f9",x"49"),
  1656 => (x"b7",x"c0",x"4b",x"70"),
  1657 => (x"fe",x"fc",x"03",x"ab"),
  1658 => (x"26",x"48",x"c0",x"87"),
  1659 => (x"26",x"4c",x"26",x"4d"),
  1660 => (x"00",x"4f",x"26",x"4b"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"1e",x"00",x"00",x"00"),
  1663 => (x"49",x"72",x"4a",x"c0"),
  1664 => (x"e9",x"c1",x"91",x"c4"),
  1665 => (x"79",x"c0",x"81",x"ca"),
  1666 => (x"b7",x"d0",x"82",x"c1"),
  1667 => (x"87",x"ee",x"04",x"aa"),
  1668 => (x"5e",x"0e",x"4f",x"26"),
  1669 => (x"0e",x"5d",x"5c",x"5b"),
  1670 => (x"e5",x"f8",x"4d",x"71"),
  1671 => (x"c4",x"4a",x"75",x"87"),
  1672 => (x"c1",x"92",x"2a",x"b7"),
  1673 => (x"75",x"82",x"ca",x"e9"),
  1674 => (x"c2",x"9c",x"cf",x"4c"),
  1675 => (x"4b",x"49",x"6a",x"94"),
  1676 => (x"9b",x"c3",x"2b",x"74"),
  1677 => (x"30",x"74",x"48",x"c2"),
  1678 => (x"bc",x"ff",x"4c",x"70"),
  1679 => (x"98",x"71",x"48",x"74"),
  1680 => (x"f5",x"f7",x"7a",x"70"),
  1681 => (x"fe",x"48",x"73",x"87"),
  1682 => (x"00",x"00",x"87",x"e1"),
  1683 => (x"00",x"00",x"00",x"00"),
  1684 => (x"00",x"00",x"00",x"00"),
  1685 => (x"00",x"00",x"00",x"00"),
  1686 => (x"00",x"00",x"00",x"00"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"00",x"00",x"00",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"00"),
  1692 => (x"00",x"00",x"00",x"00"),
  1693 => (x"00",x"00",x"00",x"00"),
  1694 => (x"00",x"00",x"00",x"00"),
  1695 => (x"00",x"00",x"00",x"00"),
  1696 => (x"00",x"00",x"00",x"00"),
  1697 => (x"00",x"00",x"00",x"00"),
  1698 => (x"ff",x"1e",x"00",x"00"),
  1699 => (x"e1",x"c8",x"48",x"d0"),
  1700 => (x"ff",x"48",x"71",x"78"),
  1701 => (x"c4",x"78",x"08",x"d4"),
  1702 => (x"d4",x"ff",x"48",x"66"),
  1703 => (x"4f",x"26",x"78",x"08"),
  1704 => (x"c4",x"4a",x"71",x"1e"),
  1705 => (x"72",x"1e",x"49",x"66"),
  1706 => (x"87",x"de",x"ff",x"49"),
  1707 => (x"c0",x"48",x"d0",x"ff"),
  1708 => (x"26",x"26",x"78",x"e0"),
  1709 => (x"1e",x"73",x"1e",x"4f"),
  1710 => (x"66",x"c8",x"4b",x"71"),
  1711 => (x"4a",x"73",x"1e",x"49"),
  1712 => (x"49",x"a2",x"e0",x"c1"),
  1713 => (x"26",x"87",x"d9",x"ff"),
  1714 => (x"4d",x"26",x"87",x"c4"),
  1715 => (x"4b",x"26",x"4c",x"26"),
  1716 => (x"ff",x"1e",x"4f",x"26"),
  1717 => (x"ff",x"c3",x"4a",x"d4"),
  1718 => (x"48",x"d0",x"ff",x"7a"),
  1719 => (x"de",x"78",x"e1",x"c0"),
  1720 => (x"d0",x"e0",x"c2",x"7a"),
  1721 => (x"48",x"49",x"7a",x"bf"),
  1722 => (x"7a",x"70",x"28",x"c8"),
  1723 => (x"28",x"d0",x"48",x"71"),
  1724 => (x"48",x"71",x"7a",x"70"),
  1725 => (x"7a",x"70",x"28",x"d8"),
  1726 => (x"c0",x"48",x"d0",x"ff"),
  1727 => (x"4f",x"26",x"78",x"e0"),
  1728 => (x"48",x"d0",x"ff",x"1e"),
  1729 => (x"71",x"78",x"c9",x"c8"),
  1730 => (x"08",x"d4",x"ff",x"48"),
  1731 => (x"1e",x"4f",x"26",x"78"),
  1732 => (x"eb",x"49",x"4a",x"71"),
  1733 => (x"48",x"d0",x"ff",x"87"),
  1734 => (x"4f",x"26",x"78",x"c8"),
  1735 => (x"71",x"1e",x"73",x"1e"),
  1736 => (x"e0",x"e0",x"c2",x"4b"),
  1737 => (x"87",x"c3",x"02",x"bf"),
  1738 => (x"ff",x"87",x"eb",x"c2"),
  1739 => (x"c9",x"c8",x"48",x"d0"),
  1740 => (x"c0",x"49",x"73",x"78"),
  1741 => (x"d4",x"ff",x"b1",x"e0"),
  1742 => (x"c2",x"78",x"71",x"48"),
  1743 => (x"c0",x"48",x"d4",x"e0"),
  1744 => (x"02",x"66",x"c8",x"78"),
  1745 => (x"ff",x"c3",x"87",x"c5"),
  1746 => (x"c0",x"87",x"c2",x"49"),
  1747 => (x"dc",x"e0",x"c2",x"49"),
  1748 => (x"02",x"66",x"cc",x"59"),
  1749 => (x"d5",x"c5",x"87",x"c6"),
  1750 => (x"87",x"c4",x"4a",x"d5"),
  1751 => (x"4a",x"ff",x"ff",x"cf"),
  1752 => (x"5a",x"e0",x"e0",x"c2"),
  1753 => (x"48",x"e0",x"e0",x"c2"),
  1754 => (x"87",x"c4",x"78",x"c1"),
  1755 => (x"4c",x"26",x"4d",x"26"),
  1756 => (x"4f",x"26",x"4b",x"26"),
  1757 => (x"5c",x"5b",x"5e",x"0e"),
  1758 => (x"4a",x"71",x"0e",x"5d"),
  1759 => (x"bf",x"dc",x"e0",x"c2"),
  1760 => (x"02",x"9a",x"72",x"4c"),
  1761 => (x"c8",x"49",x"87",x"cb"),
  1762 => (x"d2",x"ec",x"c1",x"91"),
  1763 => (x"c4",x"83",x"71",x"4b"),
  1764 => (x"d2",x"f0",x"c1",x"87"),
  1765 => (x"13",x"4d",x"c0",x"4b"),
  1766 => (x"c2",x"99",x"74",x"49"),
  1767 => (x"b9",x"bf",x"d8",x"e0"),
  1768 => (x"71",x"48",x"d4",x"ff"),
  1769 => (x"2c",x"b7",x"c1",x"78"),
  1770 => (x"ad",x"b7",x"c8",x"85"),
  1771 => (x"c2",x"87",x"e8",x"04"),
  1772 => (x"48",x"bf",x"d4",x"e0"),
  1773 => (x"e0",x"c2",x"80",x"c8"),
  1774 => (x"ef",x"fe",x"58",x"d8"),
  1775 => (x"1e",x"73",x"1e",x"87"),
  1776 => (x"4a",x"13",x"4b",x"71"),
  1777 => (x"87",x"cb",x"02",x"9a"),
  1778 => (x"e7",x"fe",x"49",x"72"),
  1779 => (x"9a",x"4a",x"13",x"87"),
  1780 => (x"fe",x"87",x"f5",x"05"),
  1781 => (x"c2",x"1e",x"87",x"da"),
  1782 => (x"49",x"bf",x"d4",x"e0"),
  1783 => (x"48",x"d4",x"e0",x"c2"),
  1784 => (x"c4",x"78",x"a1",x"c1"),
  1785 => (x"03",x"a9",x"b7",x"c0"),
  1786 => (x"d4",x"ff",x"87",x"db"),
  1787 => (x"d8",x"e0",x"c2",x"48"),
  1788 => (x"e0",x"c2",x"78",x"bf"),
  1789 => (x"c2",x"49",x"bf",x"d4"),
  1790 => (x"c1",x"48",x"d4",x"e0"),
  1791 => (x"c0",x"c4",x"78",x"a1"),
  1792 => (x"e5",x"04",x"a9",x"b7"),
  1793 => (x"48",x"d0",x"ff",x"87"),
  1794 => (x"e0",x"c2",x"78",x"c8"),
  1795 => (x"78",x"c0",x"48",x"e0"),
  1796 => (x"00",x"00",x"4f",x"26"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"5f",x"5f",x"00"),
  1800 => (x"03",x"00",x"00",x"00"),
  1801 => (x"03",x"03",x"00",x"03"),
  1802 => (x"7f",x"14",x"00",x"00"),
  1803 => (x"7f",x"7f",x"14",x"7f"),
  1804 => (x"24",x"00",x"00",x"14"),
  1805 => (x"3a",x"6b",x"6b",x"2e"),
  1806 => (x"6a",x"4c",x"00",x"12"),
  1807 => (x"56",x"6c",x"18",x"36"),
  1808 => (x"7e",x"30",x"00",x"32"),
  1809 => (x"3a",x"77",x"59",x"4f"),
  1810 => (x"00",x"00",x"40",x"68"),
  1811 => (x"00",x"03",x"07",x"04"),
  1812 => (x"00",x"00",x"00",x"00"),
  1813 => (x"41",x"63",x"3e",x"1c"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"1c",x"3e",x"63",x"41"),
  1816 => (x"2a",x"08",x"00",x"00"),
  1817 => (x"3e",x"1c",x"1c",x"3e"),
  1818 => (x"08",x"00",x"08",x"2a"),
  1819 => (x"08",x"3e",x"3e",x"08"),
  1820 => (x"00",x"00",x"00",x"08"),
  1821 => (x"00",x"60",x"e0",x"80"),
  1822 => (x"08",x"00",x"00",x"00"),
  1823 => (x"08",x"08",x"08",x"08"),
  1824 => (x"00",x"00",x"00",x"08"),
  1825 => (x"00",x"60",x"60",x"00"),
  1826 => (x"60",x"40",x"00",x"00"),
  1827 => (x"06",x"0c",x"18",x"30"),
  1828 => (x"3e",x"00",x"01",x"03"),
  1829 => (x"7f",x"4d",x"59",x"7f"),
  1830 => (x"04",x"00",x"00",x"3e"),
  1831 => (x"00",x"7f",x"7f",x"06"),
  1832 => (x"42",x"00",x"00",x"00"),
  1833 => (x"4f",x"59",x"71",x"63"),
  1834 => (x"22",x"00",x"00",x"46"),
  1835 => (x"7f",x"49",x"49",x"63"),
  1836 => (x"1c",x"18",x"00",x"36"),
  1837 => (x"7f",x"7f",x"13",x"16"),
  1838 => (x"27",x"00",x"00",x"10"),
  1839 => (x"7d",x"45",x"45",x"67"),
  1840 => (x"3c",x"00",x"00",x"39"),
  1841 => (x"79",x"49",x"4b",x"7e"),
  1842 => (x"01",x"00",x"00",x"30"),
  1843 => (x"0f",x"79",x"71",x"01"),
  1844 => (x"36",x"00",x"00",x"07"),
  1845 => (x"7f",x"49",x"49",x"7f"),
  1846 => (x"06",x"00",x"00",x"36"),
  1847 => (x"3f",x"69",x"49",x"4f"),
  1848 => (x"00",x"00",x"00",x"1e"),
  1849 => (x"00",x"66",x"66",x"00"),
  1850 => (x"00",x"00",x"00",x"00"),
  1851 => (x"00",x"66",x"e6",x"80"),
  1852 => (x"08",x"00",x"00",x"00"),
  1853 => (x"22",x"14",x"14",x"08"),
  1854 => (x"14",x"00",x"00",x"22"),
  1855 => (x"14",x"14",x"14",x"14"),
  1856 => (x"22",x"00",x"00",x"14"),
  1857 => (x"08",x"14",x"14",x"22"),
  1858 => (x"02",x"00",x"00",x"08"),
  1859 => (x"0f",x"59",x"51",x"03"),
  1860 => (x"7f",x"3e",x"00",x"06"),
  1861 => (x"1f",x"55",x"5d",x"41"),
  1862 => (x"7e",x"00",x"00",x"1e"),
  1863 => (x"7f",x"09",x"09",x"7f"),
  1864 => (x"7f",x"00",x"00",x"7e"),
  1865 => (x"7f",x"49",x"49",x"7f"),
  1866 => (x"1c",x"00",x"00",x"36"),
  1867 => (x"41",x"41",x"63",x"3e"),
  1868 => (x"7f",x"00",x"00",x"41"),
  1869 => (x"3e",x"63",x"41",x"7f"),
  1870 => (x"7f",x"00",x"00",x"1c"),
  1871 => (x"41",x"49",x"49",x"7f"),
  1872 => (x"7f",x"00",x"00",x"41"),
  1873 => (x"01",x"09",x"09",x"7f"),
  1874 => (x"3e",x"00",x"00",x"01"),
  1875 => (x"7b",x"49",x"41",x"7f"),
  1876 => (x"7f",x"00",x"00",x"7a"),
  1877 => (x"7f",x"08",x"08",x"7f"),
  1878 => (x"00",x"00",x"00",x"7f"),
  1879 => (x"41",x"7f",x"7f",x"41"),
  1880 => (x"20",x"00",x"00",x"00"),
  1881 => (x"7f",x"40",x"40",x"60"),
  1882 => (x"7f",x"7f",x"00",x"3f"),
  1883 => (x"63",x"36",x"1c",x"08"),
  1884 => (x"7f",x"00",x"00",x"41"),
  1885 => (x"40",x"40",x"40",x"7f"),
  1886 => (x"7f",x"7f",x"00",x"40"),
  1887 => (x"7f",x"06",x"0c",x"06"),
  1888 => (x"7f",x"7f",x"00",x"7f"),
  1889 => (x"7f",x"18",x"0c",x"06"),
  1890 => (x"3e",x"00",x"00",x"7f"),
  1891 => (x"7f",x"41",x"41",x"7f"),
  1892 => (x"7f",x"00",x"00",x"3e"),
  1893 => (x"0f",x"09",x"09",x"7f"),
  1894 => (x"7f",x"3e",x"00",x"06"),
  1895 => (x"7e",x"7f",x"61",x"41"),
  1896 => (x"7f",x"00",x"00",x"40"),
  1897 => (x"7f",x"19",x"09",x"7f"),
  1898 => (x"26",x"00",x"00",x"66"),
  1899 => (x"7b",x"59",x"4d",x"6f"),
  1900 => (x"01",x"00",x"00",x"32"),
  1901 => (x"01",x"7f",x"7f",x"01"),
  1902 => (x"3f",x"00",x"00",x"01"),
  1903 => (x"7f",x"40",x"40",x"7f"),
  1904 => (x"0f",x"00",x"00",x"3f"),
  1905 => (x"3f",x"70",x"70",x"3f"),
  1906 => (x"7f",x"7f",x"00",x"0f"),
  1907 => (x"7f",x"30",x"18",x"30"),
  1908 => (x"63",x"41",x"00",x"7f"),
  1909 => (x"36",x"1c",x"1c",x"36"),
  1910 => (x"03",x"01",x"41",x"63"),
  1911 => (x"06",x"7c",x"7c",x"06"),
  1912 => (x"71",x"61",x"01",x"03"),
  1913 => (x"43",x"47",x"4d",x"59"),
  1914 => (x"00",x"00",x"00",x"41"),
  1915 => (x"41",x"41",x"7f",x"7f"),
  1916 => (x"03",x"01",x"00",x"00"),
  1917 => (x"30",x"18",x"0c",x"06"),
  1918 => (x"00",x"00",x"40",x"60"),
  1919 => (x"7f",x"7f",x"41",x"41"),
  1920 => (x"0c",x"08",x"00",x"00"),
  1921 => (x"0c",x"06",x"03",x"06"),
  1922 => (x"80",x"80",x"00",x"08"),
  1923 => (x"80",x"80",x"80",x"80"),
  1924 => (x"00",x"00",x"00",x"80"),
  1925 => (x"04",x"07",x"03",x"00"),
  1926 => (x"20",x"00",x"00",x"00"),
  1927 => (x"7c",x"54",x"54",x"74"),
  1928 => (x"7f",x"00",x"00",x"78"),
  1929 => (x"7c",x"44",x"44",x"7f"),
  1930 => (x"38",x"00",x"00",x"38"),
  1931 => (x"44",x"44",x"44",x"7c"),
  1932 => (x"38",x"00",x"00",x"00"),
  1933 => (x"7f",x"44",x"44",x"7c"),
  1934 => (x"38",x"00",x"00",x"7f"),
  1935 => (x"5c",x"54",x"54",x"7c"),
  1936 => (x"04",x"00",x"00",x"18"),
  1937 => (x"05",x"05",x"7f",x"7e"),
  1938 => (x"18",x"00",x"00",x"00"),
  1939 => (x"fc",x"a4",x"a4",x"bc"),
  1940 => (x"7f",x"00",x"00",x"7c"),
  1941 => (x"7c",x"04",x"04",x"7f"),
  1942 => (x"00",x"00",x"00",x"78"),
  1943 => (x"40",x"7d",x"3d",x"00"),
  1944 => (x"80",x"00",x"00",x"00"),
  1945 => (x"7d",x"fd",x"80",x"80"),
  1946 => (x"7f",x"00",x"00",x"00"),
  1947 => (x"6c",x"38",x"10",x"7f"),
  1948 => (x"00",x"00",x"00",x"44"),
  1949 => (x"40",x"7f",x"3f",x"00"),
  1950 => (x"7c",x"7c",x"00",x"00"),
  1951 => (x"7c",x"0c",x"18",x"0c"),
  1952 => (x"7c",x"00",x"00",x"78"),
  1953 => (x"7c",x"04",x"04",x"7c"),
  1954 => (x"38",x"00",x"00",x"78"),
  1955 => (x"7c",x"44",x"44",x"7c"),
  1956 => (x"fc",x"00",x"00",x"38"),
  1957 => (x"3c",x"24",x"24",x"fc"),
  1958 => (x"18",x"00",x"00",x"18"),
  1959 => (x"fc",x"24",x"24",x"3c"),
  1960 => (x"7c",x"00",x"00",x"fc"),
  1961 => (x"0c",x"04",x"04",x"7c"),
  1962 => (x"48",x"00",x"00",x"08"),
  1963 => (x"74",x"54",x"54",x"5c"),
  1964 => (x"04",x"00",x"00",x"20"),
  1965 => (x"44",x"44",x"7f",x"3f"),
  1966 => (x"3c",x"00",x"00",x"00"),
  1967 => (x"7c",x"40",x"40",x"7c"),
  1968 => (x"1c",x"00",x"00",x"7c"),
  1969 => (x"3c",x"60",x"60",x"3c"),
  1970 => (x"7c",x"3c",x"00",x"1c"),
  1971 => (x"7c",x"60",x"30",x"60"),
  1972 => (x"6c",x"44",x"00",x"3c"),
  1973 => (x"6c",x"38",x"10",x"38"),
  1974 => (x"1c",x"00",x"00",x"44"),
  1975 => (x"3c",x"60",x"e0",x"bc"),
  1976 => (x"44",x"00",x"00",x"1c"),
  1977 => (x"4c",x"5c",x"74",x"64"),
  1978 => (x"08",x"00",x"00",x"44"),
  1979 => (x"41",x"77",x"3e",x"08"),
  1980 => (x"00",x"00",x"00",x"41"),
  1981 => (x"00",x"7f",x"7f",x"00"),
  1982 => (x"41",x"00",x"00",x"00"),
  1983 => (x"08",x"3e",x"77",x"41"),
  1984 => (x"01",x"02",x"00",x"08"),
  1985 => (x"02",x"02",x"03",x"01"),
  1986 => (x"7f",x"7f",x"00",x"01"),
  1987 => (x"7f",x"7f",x"7f",x"7f"),
  1988 => (x"08",x"08",x"00",x"7f"),
  1989 => (x"3e",x"3e",x"1c",x"1c"),
  1990 => (x"7f",x"7f",x"7f",x"7f"),
  1991 => (x"1c",x"1c",x"3e",x"3e"),
  1992 => (x"10",x"00",x"08",x"08"),
  1993 => (x"18",x"7c",x"7c",x"18"),
  1994 => (x"10",x"00",x"00",x"10"),
  1995 => (x"30",x"7c",x"7c",x"30"),
  1996 => (x"30",x"10",x"00",x"10"),
  1997 => (x"1e",x"78",x"60",x"60"),
  1998 => (x"66",x"42",x"00",x"06"),
  1999 => (x"66",x"3c",x"18",x"3c"),
  2000 => (x"38",x"78",x"00",x"42"),
  2001 => (x"6c",x"c6",x"c2",x"6a"),
  2002 => (x"00",x"60",x"00",x"38"),
  2003 => (x"00",x"00",x"60",x"00"),
  2004 => (x"5e",x"0e",x"00",x"60"),
  2005 => (x"0e",x"5d",x"5c",x"5b"),
  2006 => (x"c2",x"4c",x"71",x"1e"),
  2007 => (x"4d",x"bf",x"e5",x"e0"),
  2008 => (x"1e",x"c0",x"4b",x"c0"),
  2009 => (x"c7",x"02",x"ab",x"74"),
  2010 => (x"48",x"a6",x"c4",x"87"),
  2011 => (x"87",x"c5",x"78",x"c0"),
  2012 => (x"c1",x"48",x"a6",x"c4"),
  2013 => (x"1e",x"66",x"c4",x"78"),
  2014 => (x"df",x"ee",x"49",x"73"),
  2015 => (x"c0",x"86",x"c8",x"87"),
  2016 => (x"ef",x"ef",x"49",x"e0"),
  2017 => (x"4a",x"a5",x"c4",x"87"),
  2018 => (x"f0",x"f0",x"49",x"6a"),
  2019 => (x"87",x"c6",x"f1",x"87"),
  2020 => (x"83",x"c1",x"85",x"cb"),
  2021 => (x"04",x"ab",x"b7",x"c8"),
  2022 => (x"26",x"87",x"c7",x"ff"),
  2023 => (x"4c",x"26",x"4d",x"26"),
  2024 => (x"4f",x"26",x"4b",x"26"),
  2025 => (x"c2",x"4a",x"71",x"1e"),
  2026 => (x"c2",x"5a",x"e9",x"e0"),
  2027 => (x"c7",x"48",x"e9",x"e0"),
  2028 => (x"dd",x"fe",x"49",x"78"),
  2029 => (x"1e",x"4f",x"26",x"87"),
  2030 => (x"4a",x"71",x"1e",x"73"),
  2031 => (x"03",x"aa",x"b7",x"c0"),
  2032 => (x"ce",x"c2",x"87",x"d3"),
  2033 => (x"c4",x"05",x"bf",x"c2"),
  2034 => (x"c2",x"4b",x"c1",x"87"),
  2035 => (x"c2",x"4b",x"c0",x"87"),
  2036 => (x"c4",x"5b",x"c6",x"ce"),
  2037 => (x"c6",x"ce",x"c2",x"87"),
  2038 => (x"c2",x"ce",x"c2",x"5a"),
  2039 => (x"9a",x"c1",x"4a",x"bf"),
  2040 => (x"49",x"a2",x"c0",x"c1"),
  2041 => (x"fc",x"87",x"e8",x"ec"),
  2042 => (x"c2",x"ce",x"c2",x"48"),
  2043 => (x"ef",x"fe",x"78",x"bf"),
  2044 => (x"4a",x"71",x"1e",x"87"),
  2045 => (x"72",x"1e",x"66",x"c4"),
  2046 => (x"87",x"f9",x"ea",x"49"),
  2047 => (x"1e",x"4f",x"26",x"26"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

